module SimDualPortBRAM(
  input        clock,
  input        reset,
  input        io_wea,
  input  [7:0] io_addra,
  input  [7:0] io_addrb,
  input  [1:0] io_dina,
  output [1:0] io_douta,
  output [1:0] io_doutb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] mem_0; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_1; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_2; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_3; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_4; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_5; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_6; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_7; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_8; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_9; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_10; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_11; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_12; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_13; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_14; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_15; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_16; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_17; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_18; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_19; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_20; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_21; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_22; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_23; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_24; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_25; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_26; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_27; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_28; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_29; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_30; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_31; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_32; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_33; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_34; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_35; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_36; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_37; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_38; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_39; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_40; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_41; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_42; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_43; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_44; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_45; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_46; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_47; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_48; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_49; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_50; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_51; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_52; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_53; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_54; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_55; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_56; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_57; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_58; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_59; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_60; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_61; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_62; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_63; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_64; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_65; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_66; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_67; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_68; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_69; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_70; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_71; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_72; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_73; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_74; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_75; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_76; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_77; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_78; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_79; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_80; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_81; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_82; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_83; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_84; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_85; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_86; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_87; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_88; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_89; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_90; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_91; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_92; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_93; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_94; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_95; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_96; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_97; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_98; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_99; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_100; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_101; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_102; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_103; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_104; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_105; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_106; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_107; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_108; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_109; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_110; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_111; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_112; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_113; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_114; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_115; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_116; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_117; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_118; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_119; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_120; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_121; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_122; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_123; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_124; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_125; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_126; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_127; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_128; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_129; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_130; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_131; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_132; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_133; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_134; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_135; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_136; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_137; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_138; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_139; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_140; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_141; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_142; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_143; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_144; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_145; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_146; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_147; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_148; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_149; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_150; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_151; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_152; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_153; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_154; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_155; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_156; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_157; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_158; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_159; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_160; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_161; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_162; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_163; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_164; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_165; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_166; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_167; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_168; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_169; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_170; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_171; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_172; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_173; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_174; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_175; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_176; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_177; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_178; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_179; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_180; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_181; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_182; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_183; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_184; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_185; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_186; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_187; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_188; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_189; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_190; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_191; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_192; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_193; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_194; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_195; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_196; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_197; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_198; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_199; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_200; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_201; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_202; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_203; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_204; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_205; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_206; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_207; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_208; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_209; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_210; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_211; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_212; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_213; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_214; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_215; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_216; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_217; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_218; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_219; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_220; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_221; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_222; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_223; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_224; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_225; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_226; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_227; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_228; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_229; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_230; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_231; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_232; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_233; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_234; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_235; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_236; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_237; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_238; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_239; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_240; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_241; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_242; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_243; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_244; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_245; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_246; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_247; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_248; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_249; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_250; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_251; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_252; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_253; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_254; // @[RAMWrapper.scala 41:20]
  reg [1:0] mem_255; // @[RAMWrapper.scala 41:20]
  reg [1:0] io_douta_REG; // @[RAMWrapper.scala 43:22]
  wire [1:0] _GEN_1 = 8'h1 == io_addra ? mem_1 : mem_0; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_2 = 8'h2 == io_addra ? mem_2 : _GEN_1; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_3 = 8'h3 == io_addra ? mem_3 : _GEN_2; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_4 = 8'h4 == io_addra ? mem_4 : _GEN_3; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_5 = 8'h5 == io_addra ? mem_5 : _GEN_4; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_6 = 8'h6 == io_addra ? mem_6 : _GEN_5; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_7 = 8'h7 == io_addra ? mem_7 : _GEN_6; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_8 = 8'h8 == io_addra ? mem_8 : _GEN_7; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_9 = 8'h9 == io_addra ? mem_9 : _GEN_8; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_10 = 8'ha == io_addra ? mem_10 : _GEN_9; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_11 = 8'hb == io_addra ? mem_11 : _GEN_10; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_12 = 8'hc == io_addra ? mem_12 : _GEN_11; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_13 = 8'hd == io_addra ? mem_13 : _GEN_12; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_14 = 8'he == io_addra ? mem_14 : _GEN_13; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_15 = 8'hf == io_addra ? mem_15 : _GEN_14; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_16 = 8'h10 == io_addra ? mem_16 : _GEN_15; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_17 = 8'h11 == io_addra ? mem_17 : _GEN_16; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_18 = 8'h12 == io_addra ? mem_18 : _GEN_17; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_19 = 8'h13 == io_addra ? mem_19 : _GEN_18; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_20 = 8'h14 == io_addra ? mem_20 : _GEN_19; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_21 = 8'h15 == io_addra ? mem_21 : _GEN_20; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_22 = 8'h16 == io_addra ? mem_22 : _GEN_21; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_23 = 8'h17 == io_addra ? mem_23 : _GEN_22; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_24 = 8'h18 == io_addra ? mem_24 : _GEN_23; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_25 = 8'h19 == io_addra ? mem_25 : _GEN_24; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_26 = 8'h1a == io_addra ? mem_26 : _GEN_25; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_27 = 8'h1b == io_addra ? mem_27 : _GEN_26; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_28 = 8'h1c == io_addra ? mem_28 : _GEN_27; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_29 = 8'h1d == io_addra ? mem_29 : _GEN_28; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_30 = 8'h1e == io_addra ? mem_30 : _GEN_29; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_31 = 8'h1f == io_addra ? mem_31 : _GEN_30; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_32 = 8'h20 == io_addra ? mem_32 : _GEN_31; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_33 = 8'h21 == io_addra ? mem_33 : _GEN_32; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_34 = 8'h22 == io_addra ? mem_34 : _GEN_33; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_35 = 8'h23 == io_addra ? mem_35 : _GEN_34; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_36 = 8'h24 == io_addra ? mem_36 : _GEN_35; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_37 = 8'h25 == io_addra ? mem_37 : _GEN_36; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_38 = 8'h26 == io_addra ? mem_38 : _GEN_37; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_39 = 8'h27 == io_addra ? mem_39 : _GEN_38; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_40 = 8'h28 == io_addra ? mem_40 : _GEN_39; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_41 = 8'h29 == io_addra ? mem_41 : _GEN_40; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_42 = 8'h2a == io_addra ? mem_42 : _GEN_41; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_43 = 8'h2b == io_addra ? mem_43 : _GEN_42; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_44 = 8'h2c == io_addra ? mem_44 : _GEN_43; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_45 = 8'h2d == io_addra ? mem_45 : _GEN_44; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_46 = 8'h2e == io_addra ? mem_46 : _GEN_45; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_47 = 8'h2f == io_addra ? mem_47 : _GEN_46; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_48 = 8'h30 == io_addra ? mem_48 : _GEN_47; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_49 = 8'h31 == io_addra ? mem_49 : _GEN_48; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_50 = 8'h32 == io_addra ? mem_50 : _GEN_49; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_51 = 8'h33 == io_addra ? mem_51 : _GEN_50; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_52 = 8'h34 == io_addra ? mem_52 : _GEN_51; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_53 = 8'h35 == io_addra ? mem_53 : _GEN_52; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_54 = 8'h36 == io_addra ? mem_54 : _GEN_53; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_55 = 8'h37 == io_addra ? mem_55 : _GEN_54; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_56 = 8'h38 == io_addra ? mem_56 : _GEN_55; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_57 = 8'h39 == io_addra ? mem_57 : _GEN_56; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_58 = 8'h3a == io_addra ? mem_58 : _GEN_57; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_59 = 8'h3b == io_addra ? mem_59 : _GEN_58; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_60 = 8'h3c == io_addra ? mem_60 : _GEN_59; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_61 = 8'h3d == io_addra ? mem_61 : _GEN_60; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_62 = 8'h3e == io_addra ? mem_62 : _GEN_61; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_63 = 8'h3f == io_addra ? mem_63 : _GEN_62; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_64 = 8'h40 == io_addra ? mem_64 : _GEN_63; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_65 = 8'h41 == io_addra ? mem_65 : _GEN_64; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_66 = 8'h42 == io_addra ? mem_66 : _GEN_65; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_67 = 8'h43 == io_addra ? mem_67 : _GEN_66; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_68 = 8'h44 == io_addra ? mem_68 : _GEN_67; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_69 = 8'h45 == io_addra ? mem_69 : _GEN_68; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_70 = 8'h46 == io_addra ? mem_70 : _GEN_69; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_71 = 8'h47 == io_addra ? mem_71 : _GEN_70; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_72 = 8'h48 == io_addra ? mem_72 : _GEN_71; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_73 = 8'h49 == io_addra ? mem_73 : _GEN_72; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_74 = 8'h4a == io_addra ? mem_74 : _GEN_73; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_75 = 8'h4b == io_addra ? mem_75 : _GEN_74; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_76 = 8'h4c == io_addra ? mem_76 : _GEN_75; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_77 = 8'h4d == io_addra ? mem_77 : _GEN_76; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_78 = 8'h4e == io_addra ? mem_78 : _GEN_77; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_79 = 8'h4f == io_addra ? mem_79 : _GEN_78; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_80 = 8'h50 == io_addra ? mem_80 : _GEN_79; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_81 = 8'h51 == io_addra ? mem_81 : _GEN_80; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_82 = 8'h52 == io_addra ? mem_82 : _GEN_81; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_83 = 8'h53 == io_addra ? mem_83 : _GEN_82; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_84 = 8'h54 == io_addra ? mem_84 : _GEN_83; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_85 = 8'h55 == io_addra ? mem_85 : _GEN_84; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_86 = 8'h56 == io_addra ? mem_86 : _GEN_85; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_87 = 8'h57 == io_addra ? mem_87 : _GEN_86; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_88 = 8'h58 == io_addra ? mem_88 : _GEN_87; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_89 = 8'h59 == io_addra ? mem_89 : _GEN_88; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_90 = 8'h5a == io_addra ? mem_90 : _GEN_89; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_91 = 8'h5b == io_addra ? mem_91 : _GEN_90; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_92 = 8'h5c == io_addra ? mem_92 : _GEN_91; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_93 = 8'h5d == io_addra ? mem_93 : _GEN_92; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_94 = 8'h5e == io_addra ? mem_94 : _GEN_93; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_95 = 8'h5f == io_addra ? mem_95 : _GEN_94; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_96 = 8'h60 == io_addra ? mem_96 : _GEN_95; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_97 = 8'h61 == io_addra ? mem_97 : _GEN_96; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_98 = 8'h62 == io_addra ? mem_98 : _GEN_97; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_99 = 8'h63 == io_addra ? mem_99 : _GEN_98; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_100 = 8'h64 == io_addra ? mem_100 : _GEN_99; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_101 = 8'h65 == io_addra ? mem_101 : _GEN_100; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_102 = 8'h66 == io_addra ? mem_102 : _GEN_101; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_103 = 8'h67 == io_addra ? mem_103 : _GEN_102; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_104 = 8'h68 == io_addra ? mem_104 : _GEN_103; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_105 = 8'h69 == io_addra ? mem_105 : _GEN_104; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_106 = 8'h6a == io_addra ? mem_106 : _GEN_105; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_107 = 8'h6b == io_addra ? mem_107 : _GEN_106; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_108 = 8'h6c == io_addra ? mem_108 : _GEN_107; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_109 = 8'h6d == io_addra ? mem_109 : _GEN_108; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_110 = 8'h6e == io_addra ? mem_110 : _GEN_109; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_111 = 8'h6f == io_addra ? mem_111 : _GEN_110; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_112 = 8'h70 == io_addra ? mem_112 : _GEN_111; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_113 = 8'h71 == io_addra ? mem_113 : _GEN_112; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_114 = 8'h72 == io_addra ? mem_114 : _GEN_113; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_115 = 8'h73 == io_addra ? mem_115 : _GEN_114; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_116 = 8'h74 == io_addra ? mem_116 : _GEN_115; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_117 = 8'h75 == io_addra ? mem_117 : _GEN_116; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_118 = 8'h76 == io_addra ? mem_118 : _GEN_117; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_119 = 8'h77 == io_addra ? mem_119 : _GEN_118; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_120 = 8'h78 == io_addra ? mem_120 : _GEN_119; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_121 = 8'h79 == io_addra ? mem_121 : _GEN_120; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_122 = 8'h7a == io_addra ? mem_122 : _GEN_121; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_123 = 8'h7b == io_addra ? mem_123 : _GEN_122; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_124 = 8'h7c == io_addra ? mem_124 : _GEN_123; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_125 = 8'h7d == io_addra ? mem_125 : _GEN_124; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_126 = 8'h7e == io_addra ? mem_126 : _GEN_125; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_127 = 8'h7f == io_addra ? mem_127 : _GEN_126; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_128 = 8'h80 == io_addra ? mem_128 : _GEN_127; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_129 = 8'h81 == io_addra ? mem_129 : _GEN_128; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_130 = 8'h82 == io_addra ? mem_130 : _GEN_129; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_131 = 8'h83 == io_addra ? mem_131 : _GEN_130; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_132 = 8'h84 == io_addra ? mem_132 : _GEN_131; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_133 = 8'h85 == io_addra ? mem_133 : _GEN_132; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_134 = 8'h86 == io_addra ? mem_134 : _GEN_133; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_135 = 8'h87 == io_addra ? mem_135 : _GEN_134; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_136 = 8'h88 == io_addra ? mem_136 : _GEN_135; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_137 = 8'h89 == io_addra ? mem_137 : _GEN_136; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_138 = 8'h8a == io_addra ? mem_138 : _GEN_137; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_139 = 8'h8b == io_addra ? mem_139 : _GEN_138; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_140 = 8'h8c == io_addra ? mem_140 : _GEN_139; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_141 = 8'h8d == io_addra ? mem_141 : _GEN_140; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_142 = 8'h8e == io_addra ? mem_142 : _GEN_141; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_143 = 8'h8f == io_addra ? mem_143 : _GEN_142; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_144 = 8'h90 == io_addra ? mem_144 : _GEN_143; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_145 = 8'h91 == io_addra ? mem_145 : _GEN_144; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_146 = 8'h92 == io_addra ? mem_146 : _GEN_145; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_147 = 8'h93 == io_addra ? mem_147 : _GEN_146; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_148 = 8'h94 == io_addra ? mem_148 : _GEN_147; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_149 = 8'h95 == io_addra ? mem_149 : _GEN_148; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_150 = 8'h96 == io_addra ? mem_150 : _GEN_149; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_151 = 8'h97 == io_addra ? mem_151 : _GEN_150; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_152 = 8'h98 == io_addra ? mem_152 : _GEN_151; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_153 = 8'h99 == io_addra ? mem_153 : _GEN_152; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_154 = 8'h9a == io_addra ? mem_154 : _GEN_153; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_155 = 8'h9b == io_addra ? mem_155 : _GEN_154; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_156 = 8'h9c == io_addra ? mem_156 : _GEN_155; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_157 = 8'h9d == io_addra ? mem_157 : _GEN_156; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_158 = 8'h9e == io_addra ? mem_158 : _GEN_157; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_159 = 8'h9f == io_addra ? mem_159 : _GEN_158; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_160 = 8'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_161 = 8'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_162 = 8'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_163 = 8'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_164 = 8'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_165 = 8'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_166 = 8'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_167 = 8'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_168 = 8'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_169 = 8'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_170 = 8'haa == io_addra ? mem_170 : _GEN_169; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_171 = 8'hab == io_addra ? mem_171 : _GEN_170; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_172 = 8'hac == io_addra ? mem_172 : _GEN_171; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_173 = 8'had == io_addra ? mem_173 : _GEN_172; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_174 = 8'hae == io_addra ? mem_174 : _GEN_173; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_175 = 8'haf == io_addra ? mem_175 : _GEN_174; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_176 = 8'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_177 = 8'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_178 = 8'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_179 = 8'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_180 = 8'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_181 = 8'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_182 = 8'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_183 = 8'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_184 = 8'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_185 = 8'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_186 = 8'hba == io_addra ? mem_186 : _GEN_185; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_187 = 8'hbb == io_addra ? mem_187 : _GEN_186; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_188 = 8'hbc == io_addra ? mem_188 : _GEN_187; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_189 = 8'hbd == io_addra ? mem_189 : _GEN_188; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_190 = 8'hbe == io_addra ? mem_190 : _GEN_189; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_191 = 8'hbf == io_addra ? mem_191 : _GEN_190; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_192 = 8'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_193 = 8'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_194 = 8'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_195 = 8'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_196 = 8'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_197 = 8'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_198 = 8'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_199 = 8'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_200 = 8'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_201 = 8'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_202 = 8'hca == io_addra ? mem_202 : _GEN_201; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_203 = 8'hcb == io_addra ? mem_203 : _GEN_202; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_204 = 8'hcc == io_addra ? mem_204 : _GEN_203; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_205 = 8'hcd == io_addra ? mem_205 : _GEN_204; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_206 = 8'hce == io_addra ? mem_206 : _GEN_205; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_207 = 8'hcf == io_addra ? mem_207 : _GEN_206; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_208 = 8'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_209 = 8'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_210 = 8'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_211 = 8'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_212 = 8'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_213 = 8'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_214 = 8'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_215 = 8'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_216 = 8'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_217 = 8'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_218 = 8'hda == io_addra ? mem_218 : _GEN_217; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_219 = 8'hdb == io_addra ? mem_219 : _GEN_218; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_220 = 8'hdc == io_addra ? mem_220 : _GEN_219; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_221 = 8'hdd == io_addra ? mem_221 : _GEN_220; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_222 = 8'hde == io_addra ? mem_222 : _GEN_221; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_223 = 8'hdf == io_addra ? mem_223 : _GEN_222; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_224 = 8'he0 == io_addra ? mem_224 : _GEN_223; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_225 = 8'he1 == io_addra ? mem_225 : _GEN_224; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_226 = 8'he2 == io_addra ? mem_226 : _GEN_225; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_227 = 8'he3 == io_addra ? mem_227 : _GEN_226; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_228 = 8'he4 == io_addra ? mem_228 : _GEN_227; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_229 = 8'he5 == io_addra ? mem_229 : _GEN_228; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_230 = 8'he6 == io_addra ? mem_230 : _GEN_229; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_231 = 8'he7 == io_addra ? mem_231 : _GEN_230; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_232 = 8'he8 == io_addra ? mem_232 : _GEN_231; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_233 = 8'he9 == io_addra ? mem_233 : _GEN_232; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_234 = 8'hea == io_addra ? mem_234 : _GEN_233; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_235 = 8'heb == io_addra ? mem_235 : _GEN_234; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_236 = 8'hec == io_addra ? mem_236 : _GEN_235; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_237 = 8'hed == io_addra ? mem_237 : _GEN_236; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_238 = 8'hee == io_addra ? mem_238 : _GEN_237; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_239 = 8'hef == io_addra ? mem_239 : _GEN_238; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_240 = 8'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_241 = 8'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_242 = 8'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_243 = 8'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_244 = 8'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_245 = 8'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_246 = 8'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_247 = 8'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_248 = 8'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_249 = 8'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_250 = 8'hfa == io_addra ? mem_250 : _GEN_249; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [1:0] _GEN_251 = 8'hfb == io_addra ? mem_251 : _GEN_250; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  reg [1:0] io_doutb_REG; // @[RAMWrapper.scala 44:22]
  wire [1:0] _GEN_257 = 8'h1 == io_addrb ? mem_1 : mem_0; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_258 = 8'h2 == io_addrb ? mem_2 : _GEN_257; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_259 = 8'h3 == io_addrb ? mem_3 : _GEN_258; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_260 = 8'h4 == io_addrb ? mem_4 : _GEN_259; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_261 = 8'h5 == io_addrb ? mem_5 : _GEN_260; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_262 = 8'h6 == io_addrb ? mem_6 : _GEN_261; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_263 = 8'h7 == io_addrb ? mem_7 : _GEN_262; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_264 = 8'h8 == io_addrb ? mem_8 : _GEN_263; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_265 = 8'h9 == io_addrb ? mem_9 : _GEN_264; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_266 = 8'ha == io_addrb ? mem_10 : _GEN_265; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_267 = 8'hb == io_addrb ? mem_11 : _GEN_266; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_268 = 8'hc == io_addrb ? mem_12 : _GEN_267; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_269 = 8'hd == io_addrb ? mem_13 : _GEN_268; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_270 = 8'he == io_addrb ? mem_14 : _GEN_269; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_271 = 8'hf == io_addrb ? mem_15 : _GEN_270; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_272 = 8'h10 == io_addrb ? mem_16 : _GEN_271; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_273 = 8'h11 == io_addrb ? mem_17 : _GEN_272; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_274 = 8'h12 == io_addrb ? mem_18 : _GEN_273; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_275 = 8'h13 == io_addrb ? mem_19 : _GEN_274; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_276 = 8'h14 == io_addrb ? mem_20 : _GEN_275; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_277 = 8'h15 == io_addrb ? mem_21 : _GEN_276; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_278 = 8'h16 == io_addrb ? mem_22 : _GEN_277; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_279 = 8'h17 == io_addrb ? mem_23 : _GEN_278; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_280 = 8'h18 == io_addrb ? mem_24 : _GEN_279; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_281 = 8'h19 == io_addrb ? mem_25 : _GEN_280; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_282 = 8'h1a == io_addrb ? mem_26 : _GEN_281; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_283 = 8'h1b == io_addrb ? mem_27 : _GEN_282; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_284 = 8'h1c == io_addrb ? mem_28 : _GEN_283; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_285 = 8'h1d == io_addrb ? mem_29 : _GEN_284; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_286 = 8'h1e == io_addrb ? mem_30 : _GEN_285; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_287 = 8'h1f == io_addrb ? mem_31 : _GEN_286; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_288 = 8'h20 == io_addrb ? mem_32 : _GEN_287; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_289 = 8'h21 == io_addrb ? mem_33 : _GEN_288; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_290 = 8'h22 == io_addrb ? mem_34 : _GEN_289; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_291 = 8'h23 == io_addrb ? mem_35 : _GEN_290; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_292 = 8'h24 == io_addrb ? mem_36 : _GEN_291; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_293 = 8'h25 == io_addrb ? mem_37 : _GEN_292; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_294 = 8'h26 == io_addrb ? mem_38 : _GEN_293; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_295 = 8'h27 == io_addrb ? mem_39 : _GEN_294; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_296 = 8'h28 == io_addrb ? mem_40 : _GEN_295; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_297 = 8'h29 == io_addrb ? mem_41 : _GEN_296; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_298 = 8'h2a == io_addrb ? mem_42 : _GEN_297; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_299 = 8'h2b == io_addrb ? mem_43 : _GEN_298; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_300 = 8'h2c == io_addrb ? mem_44 : _GEN_299; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_301 = 8'h2d == io_addrb ? mem_45 : _GEN_300; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_302 = 8'h2e == io_addrb ? mem_46 : _GEN_301; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_303 = 8'h2f == io_addrb ? mem_47 : _GEN_302; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_304 = 8'h30 == io_addrb ? mem_48 : _GEN_303; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_305 = 8'h31 == io_addrb ? mem_49 : _GEN_304; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_306 = 8'h32 == io_addrb ? mem_50 : _GEN_305; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_307 = 8'h33 == io_addrb ? mem_51 : _GEN_306; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_308 = 8'h34 == io_addrb ? mem_52 : _GEN_307; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_309 = 8'h35 == io_addrb ? mem_53 : _GEN_308; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_310 = 8'h36 == io_addrb ? mem_54 : _GEN_309; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_311 = 8'h37 == io_addrb ? mem_55 : _GEN_310; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_312 = 8'h38 == io_addrb ? mem_56 : _GEN_311; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_313 = 8'h39 == io_addrb ? mem_57 : _GEN_312; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_314 = 8'h3a == io_addrb ? mem_58 : _GEN_313; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_315 = 8'h3b == io_addrb ? mem_59 : _GEN_314; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_316 = 8'h3c == io_addrb ? mem_60 : _GEN_315; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_317 = 8'h3d == io_addrb ? mem_61 : _GEN_316; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_318 = 8'h3e == io_addrb ? mem_62 : _GEN_317; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_319 = 8'h3f == io_addrb ? mem_63 : _GEN_318; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_320 = 8'h40 == io_addrb ? mem_64 : _GEN_319; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_321 = 8'h41 == io_addrb ? mem_65 : _GEN_320; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_322 = 8'h42 == io_addrb ? mem_66 : _GEN_321; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_323 = 8'h43 == io_addrb ? mem_67 : _GEN_322; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_324 = 8'h44 == io_addrb ? mem_68 : _GEN_323; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_325 = 8'h45 == io_addrb ? mem_69 : _GEN_324; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_326 = 8'h46 == io_addrb ? mem_70 : _GEN_325; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_327 = 8'h47 == io_addrb ? mem_71 : _GEN_326; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_328 = 8'h48 == io_addrb ? mem_72 : _GEN_327; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_329 = 8'h49 == io_addrb ? mem_73 : _GEN_328; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_330 = 8'h4a == io_addrb ? mem_74 : _GEN_329; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_331 = 8'h4b == io_addrb ? mem_75 : _GEN_330; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_332 = 8'h4c == io_addrb ? mem_76 : _GEN_331; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_333 = 8'h4d == io_addrb ? mem_77 : _GEN_332; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_334 = 8'h4e == io_addrb ? mem_78 : _GEN_333; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_335 = 8'h4f == io_addrb ? mem_79 : _GEN_334; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_336 = 8'h50 == io_addrb ? mem_80 : _GEN_335; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_337 = 8'h51 == io_addrb ? mem_81 : _GEN_336; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_338 = 8'h52 == io_addrb ? mem_82 : _GEN_337; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_339 = 8'h53 == io_addrb ? mem_83 : _GEN_338; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_340 = 8'h54 == io_addrb ? mem_84 : _GEN_339; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_341 = 8'h55 == io_addrb ? mem_85 : _GEN_340; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_342 = 8'h56 == io_addrb ? mem_86 : _GEN_341; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_343 = 8'h57 == io_addrb ? mem_87 : _GEN_342; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_344 = 8'h58 == io_addrb ? mem_88 : _GEN_343; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_345 = 8'h59 == io_addrb ? mem_89 : _GEN_344; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_346 = 8'h5a == io_addrb ? mem_90 : _GEN_345; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_347 = 8'h5b == io_addrb ? mem_91 : _GEN_346; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_348 = 8'h5c == io_addrb ? mem_92 : _GEN_347; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_349 = 8'h5d == io_addrb ? mem_93 : _GEN_348; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_350 = 8'h5e == io_addrb ? mem_94 : _GEN_349; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_351 = 8'h5f == io_addrb ? mem_95 : _GEN_350; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_352 = 8'h60 == io_addrb ? mem_96 : _GEN_351; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_353 = 8'h61 == io_addrb ? mem_97 : _GEN_352; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_354 = 8'h62 == io_addrb ? mem_98 : _GEN_353; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_355 = 8'h63 == io_addrb ? mem_99 : _GEN_354; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_356 = 8'h64 == io_addrb ? mem_100 : _GEN_355; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_357 = 8'h65 == io_addrb ? mem_101 : _GEN_356; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_358 = 8'h66 == io_addrb ? mem_102 : _GEN_357; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_359 = 8'h67 == io_addrb ? mem_103 : _GEN_358; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_360 = 8'h68 == io_addrb ? mem_104 : _GEN_359; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_361 = 8'h69 == io_addrb ? mem_105 : _GEN_360; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_362 = 8'h6a == io_addrb ? mem_106 : _GEN_361; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_363 = 8'h6b == io_addrb ? mem_107 : _GEN_362; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_364 = 8'h6c == io_addrb ? mem_108 : _GEN_363; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_365 = 8'h6d == io_addrb ? mem_109 : _GEN_364; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_366 = 8'h6e == io_addrb ? mem_110 : _GEN_365; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_367 = 8'h6f == io_addrb ? mem_111 : _GEN_366; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_368 = 8'h70 == io_addrb ? mem_112 : _GEN_367; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_369 = 8'h71 == io_addrb ? mem_113 : _GEN_368; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_370 = 8'h72 == io_addrb ? mem_114 : _GEN_369; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_371 = 8'h73 == io_addrb ? mem_115 : _GEN_370; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_372 = 8'h74 == io_addrb ? mem_116 : _GEN_371; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_373 = 8'h75 == io_addrb ? mem_117 : _GEN_372; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_374 = 8'h76 == io_addrb ? mem_118 : _GEN_373; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_375 = 8'h77 == io_addrb ? mem_119 : _GEN_374; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_376 = 8'h78 == io_addrb ? mem_120 : _GEN_375; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_377 = 8'h79 == io_addrb ? mem_121 : _GEN_376; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_378 = 8'h7a == io_addrb ? mem_122 : _GEN_377; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_379 = 8'h7b == io_addrb ? mem_123 : _GEN_378; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_380 = 8'h7c == io_addrb ? mem_124 : _GEN_379; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_381 = 8'h7d == io_addrb ? mem_125 : _GEN_380; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_382 = 8'h7e == io_addrb ? mem_126 : _GEN_381; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_383 = 8'h7f == io_addrb ? mem_127 : _GEN_382; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_384 = 8'h80 == io_addrb ? mem_128 : _GEN_383; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_385 = 8'h81 == io_addrb ? mem_129 : _GEN_384; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_386 = 8'h82 == io_addrb ? mem_130 : _GEN_385; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_387 = 8'h83 == io_addrb ? mem_131 : _GEN_386; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_388 = 8'h84 == io_addrb ? mem_132 : _GEN_387; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_389 = 8'h85 == io_addrb ? mem_133 : _GEN_388; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_390 = 8'h86 == io_addrb ? mem_134 : _GEN_389; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_391 = 8'h87 == io_addrb ? mem_135 : _GEN_390; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_392 = 8'h88 == io_addrb ? mem_136 : _GEN_391; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_393 = 8'h89 == io_addrb ? mem_137 : _GEN_392; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_394 = 8'h8a == io_addrb ? mem_138 : _GEN_393; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_395 = 8'h8b == io_addrb ? mem_139 : _GEN_394; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_396 = 8'h8c == io_addrb ? mem_140 : _GEN_395; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_397 = 8'h8d == io_addrb ? mem_141 : _GEN_396; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_398 = 8'h8e == io_addrb ? mem_142 : _GEN_397; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_399 = 8'h8f == io_addrb ? mem_143 : _GEN_398; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_400 = 8'h90 == io_addrb ? mem_144 : _GEN_399; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_401 = 8'h91 == io_addrb ? mem_145 : _GEN_400; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_402 = 8'h92 == io_addrb ? mem_146 : _GEN_401; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_403 = 8'h93 == io_addrb ? mem_147 : _GEN_402; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_404 = 8'h94 == io_addrb ? mem_148 : _GEN_403; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_405 = 8'h95 == io_addrb ? mem_149 : _GEN_404; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_406 = 8'h96 == io_addrb ? mem_150 : _GEN_405; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_407 = 8'h97 == io_addrb ? mem_151 : _GEN_406; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_408 = 8'h98 == io_addrb ? mem_152 : _GEN_407; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_409 = 8'h99 == io_addrb ? mem_153 : _GEN_408; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_410 = 8'h9a == io_addrb ? mem_154 : _GEN_409; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_411 = 8'h9b == io_addrb ? mem_155 : _GEN_410; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_412 = 8'h9c == io_addrb ? mem_156 : _GEN_411; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_413 = 8'h9d == io_addrb ? mem_157 : _GEN_412; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_414 = 8'h9e == io_addrb ? mem_158 : _GEN_413; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_415 = 8'h9f == io_addrb ? mem_159 : _GEN_414; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_416 = 8'ha0 == io_addrb ? mem_160 : _GEN_415; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_417 = 8'ha1 == io_addrb ? mem_161 : _GEN_416; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_418 = 8'ha2 == io_addrb ? mem_162 : _GEN_417; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_419 = 8'ha3 == io_addrb ? mem_163 : _GEN_418; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_420 = 8'ha4 == io_addrb ? mem_164 : _GEN_419; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_421 = 8'ha5 == io_addrb ? mem_165 : _GEN_420; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_422 = 8'ha6 == io_addrb ? mem_166 : _GEN_421; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_423 = 8'ha7 == io_addrb ? mem_167 : _GEN_422; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_424 = 8'ha8 == io_addrb ? mem_168 : _GEN_423; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_425 = 8'ha9 == io_addrb ? mem_169 : _GEN_424; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_426 = 8'haa == io_addrb ? mem_170 : _GEN_425; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_427 = 8'hab == io_addrb ? mem_171 : _GEN_426; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_428 = 8'hac == io_addrb ? mem_172 : _GEN_427; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_429 = 8'had == io_addrb ? mem_173 : _GEN_428; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_430 = 8'hae == io_addrb ? mem_174 : _GEN_429; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_431 = 8'haf == io_addrb ? mem_175 : _GEN_430; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_432 = 8'hb0 == io_addrb ? mem_176 : _GEN_431; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_433 = 8'hb1 == io_addrb ? mem_177 : _GEN_432; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_434 = 8'hb2 == io_addrb ? mem_178 : _GEN_433; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_435 = 8'hb3 == io_addrb ? mem_179 : _GEN_434; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_436 = 8'hb4 == io_addrb ? mem_180 : _GEN_435; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_437 = 8'hb5 == io_addrb ? mem_181 : _GEN_436; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_438 = 8'hb6 == io_addrb ? mem_182 : _GEN_437; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_439 = 8'hb7 == io_addrb ? mem_183 : _GEN_438; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_440 = 8'hb8 == io_addrb ? mem_184 : _GEN_439; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_441 = 8'hb9 == io_addrb ? mem_185 : _GEN_440; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_442 = 8'hba == io_addrb ? mem_186 : _GEN_441; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_443 = 8'hbb == io_addrb ? mem_187 : _GEN_442; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_444 = 8'hbc == io_addrb ? mem_188 : _GEN_443; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_445 = 8'hbd == io_addrb ? mem_189 : _GEN_444; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_446 = 8'hbe == io_addrb ? mem_190 : _GEN_445; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_447 = 8'hbf == io_addrb ? mem_191 : _GEN_446; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_448 = 8'hc0 == io_addrb ? mem_192 : _GEN_447; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_449 = 8'hc1 == io_addrb ? mem_193 : _GEN_448; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_450 = 8'hc2 == io_addrb ? mem_194 : _GEN_449; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_451 = 8'hc3 == io_addrb ? mem_195 : _GEN_450; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_452 = 8'hc4 == io_addrb ? mem_196 : _GEN_451; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_453 = 8'hc5 == io_addrb ? mem_197 : _GEN_452; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_454 = 8'hc6 == io_addrb ? mem_198 : _GEN_453; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_455 = 8'hc7 == io_addrb ? mem_199 : _GEN_454; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_456 = 8'hc8 == io_addrb ? mem_200 : _GEN_455; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_457 = 8'hc9 == io_addrb ? mem_201 : _GEN_456; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_458 = 8'hca == io_addrb ? mem_202 : _GEN_457; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_459 = 8'hcb == io_addrb ? mem_203 : _GEN_458; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_460 = 8'hcc == io_addrb ? mem_204 : _GEN_459; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_461 = 8'hcd == io_addrb ? mem_205 : _GEN_460; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_462 = 8'hce == io_addrb ? mem_206 : _GEN_461; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_463 = 8'hcf == io_addrb ? mem_207 : _GEN_462; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_464 = 8'hd0 == io_addrb ? mem_208 : _GEN_463; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_465 = 8'hd1 == io_addrb ? mem_209 : _GEN_464; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_466 = 8'hd2 == io_addrb ? mem_210 : _GEN_465; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_467 = 8'hd3 == io_addrb ? mem_211 : _GEN_466; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_468 = 8'hd4 == io_addrb ? mem_212 : _GEN_467; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_469 = 8'hd5 == io_addrb ? mem_213 : _GEN_468; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_470 = 8'hd6 == io_addrb ? mem_214 : _GEN_469; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_471 = 8'hd7 == io_addrb ? mem_215 : _GEN_470; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_472 = 8'hd8 == io_addrb ? mem_216 : _GEN_471; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_473 = 8'hd9 == io_addrb ? mem_217 : _GEN_472; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_474 = 8'hda == io_addrb ? mem_218 : _GEN_473; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_475 = 8'hdb == io_addrb ? mem_219 : _GEN_474; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_476 = 8'hdc == io_addrb ? mem_220 : _GEN_475; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_477 = 8'hdd == io_addrb ? mem_221 : _GEN_476; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_478 = 8'hde == io_addrb ? mem_222 : _GEN_477; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_479 = 8'hdf == io_addrb ? mem_223 : _GEN_478; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_480 = 8'he0 == io_addrb ? mem_224 : _GEN_479; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_481 = 8'he1 == io_addrb ? mem_225 : _GEN_480; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_482 = 8'he2 == io_addrb ? mem_226 : _GEN_481; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_483 = 8'he3 == io_addrb ? mem_227 : _GEN_482; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_484 = 8'he4 == io_addrb ? mem_228 : _GEN_483; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_485 = 8'he5 == io_addrb ? mem_229 : _GEN_484; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_486 = 8'he6 == io_addrb ? mem_230 : _GEN_485; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_487 = 8'he7 == io_addrb ? mem_231 : _GEN_486; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_488 = 8'he8 == io_addrb ? mem_232 : _GEN_487; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_489 = 8'he9 == io_addrb ? mem_233 : _GEN_488; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_490 = 8'hea == io_addrb ? mem_234 : _GEN_489; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_491 = 8'heb == io_addrb ? mem_235 : _GEN_490; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_492 = 8'hec == io_addrb ? mem_236 : _GEN_491; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_493 = 8'hed == io_addrb ? mem_237 : _GEN_492; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_494 = 8'hee == io_addrb ? mem_238 : _GEN_493; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_495 = 8'hef == io_addrb ? mem_239 : _GEN_494; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_496 = 8'hf0 == io_addrb ? mem_240 : _GEN_495; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_497 = 8'hf1 == io_addrb ? mem_241 : _GEN_496; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_498 = 8'hf2 == io_addrb ? mem_242 : _GEN_497; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_499 = 8'hf3 == io_addrb ? mem_243 : _GEN_498; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_500 = 8'hf4 == io_addrb ? mem_244 : _GEN_499; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_501 = 8'hf5 == io_addrb ? mem_245 : _GEN_500; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_502 = 8'hf6 == io_addrb ? mem_246 : _GEN_501; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_503 = 8'hf7 == io_addrb ? mem_247 : _GEN_502; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_504 = 8'hf8 == io_addrb ? mem_248 : _GEN_503; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_505 = 8'hf9 == io_addrb ? mem_249 : _GEN_504; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_506 = 8'hfa == io_addrb ? mem_250 : _GEN_505; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [1:0] _GEN_507 = 8'hfb == io_addrb ? mem_251 : _GEN_506; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  assign io_douta = io_douta_REG; // @[RAMWrapper.scala 43:12]
  assign io_doutb = io_doutb_REG; // @[RAMWrapper.scala 44:12]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_0 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_0 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_1 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_1 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_2 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_2 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_3 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_3 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_4 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_4 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_5 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_5 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_6 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_6 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_7 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_7 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_8 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_8 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_9 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_9 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_10 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_10 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_11 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_11 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_12 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_12 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_13 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_13 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_14 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_14 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_15 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_15 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_16 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h10 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_16 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_17 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h11 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_17 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_18 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h12 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_18 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_19 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h13 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_19 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_20 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h14 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_20 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_21 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h15 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_21 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_22 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h16 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_22 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_23 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h17 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_23 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_24 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h18 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_24 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_25 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h19 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_25 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_26 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_26 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_27 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_27 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_28 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_28 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_29 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_29 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_30 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_30 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_31 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_31 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_32 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h20 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_32 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_33 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h21 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_33 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_34 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h22 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_34 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_35 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h23 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_35 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_36 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h24 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_36 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_37 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h25 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_37 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_38 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h26 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_38 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_39 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h27 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_39 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_40 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h28 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_40 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_41 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h29 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_41 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_42 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_42 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_43 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_43 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_44 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_44 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_45 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_45 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_46 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_46 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_47 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_47 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_48 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h30 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_48 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_49 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h31 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_49 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_50 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h32 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_50 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_51 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h33 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_51 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_52 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h34 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_52 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_53 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h35 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_53 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_54 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h36 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_54 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_55 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h37 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_55 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_56 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h38 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_56 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_57 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h39 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_57 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_58 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_58 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_59 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_59 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_60 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_60 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_61 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_61 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_62 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_62 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_63 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_63 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_64 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h40 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_64 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_65 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h41 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_65 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_66 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h42 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_66 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_67 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h43 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_67 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_68 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h44 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_68 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_69 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h45 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_69 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_70 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h46 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_70 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_71 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h47 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_71 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_72 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h48 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_72 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_73 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h49 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_73 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_74 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_74 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_75 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_75 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_76 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_76 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_77 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_77 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_78 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_78 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_79 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_79 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_80 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h50 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_80 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_81 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h51 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_81 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_82 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h52 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_82 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_83 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h53 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_83 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_84 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h54 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_84 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_85 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h55 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_85 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_86 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h56 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_86 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_87 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h57 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_87 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_88 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h58 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_88 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_89 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h59 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_89 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_90 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_90 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_91 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_91 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_92 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_92 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_93 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_93 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_94 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_94 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_95 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_95 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_96 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h60 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_96 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_97 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h61 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_97 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_98 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h62 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_98 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_99 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h63 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_99 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_100 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h64 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_100 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_101 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h65 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_101 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_102 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h66 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_102 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_103 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h67 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_103 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_104 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h68 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_104 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_105 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h69 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_105 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_106 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_106 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_107 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_107 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_108 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_108 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_109 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_109 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_110 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_110 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_111 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_111 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_112 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h70 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_112 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_113 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h71 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_113 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_114 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h72 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_114 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_115 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h73 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_115 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_116 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h74 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_116 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_117 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h75 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_117 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_118 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h76 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_118 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_119 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h77 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_119 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_120 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h78 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_120 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_121 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h79 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_121 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_122 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_122 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_123 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_123 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_124 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_124 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_125 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_125 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_126 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_126 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_127 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_127 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_128 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h80 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_128 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_129 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h81 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_129 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_130 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h82 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_130 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_131 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h83 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_131 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_132 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h84 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_132 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_133 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h85 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_133 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_134 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h86 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_134 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_135 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h87 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_135 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_136 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h88 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_136 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_137 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h89 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_137 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_138 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_138 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_139 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_139 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_140 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_140 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_141 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_141 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_142 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_142 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_143 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_143 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_144 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h90 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_144 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_145 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h91 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_145 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_146 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h92 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_146 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_147 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h93 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_147 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_148 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h94 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_148 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_149 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h95 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_149 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_150 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h96 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_150 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_151 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h97 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_151 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_152 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h98 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_152 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_153 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h99 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_153 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_154 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_154 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_155 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_155 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_156 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_156 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_157 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_157 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_158 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_158 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_159 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_159 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_160 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_160 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_161 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_161 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_162 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_162 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_163 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_163 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_164 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_164 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_165 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_165 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_166 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_166 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_167 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_167 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_168 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_168 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_169 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_169 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_170 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'haa == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_170 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_171 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hab == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_171 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_172 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hac == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_172 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_173 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'had == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_173 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_174 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hae == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_174 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_175 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'haf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_175 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_176 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_176 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_177 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_177 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_178 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_178 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_179 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_179 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_180 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_180 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_181 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_181 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_182 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_182 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_183 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_183 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_184 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_184 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_185 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_185 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_186 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hba == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_186 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_187 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_187 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_188 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_188 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_189 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_189 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_190 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbe == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_190 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_191 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_191 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_192 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_192 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_193 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_193 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_194 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_194 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_195 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_195 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_196 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_196 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_197 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_197 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_198 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_198 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_199 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_199 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_200 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_200 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_201 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_201 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_202 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hca == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_202 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_203 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_203 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_204 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_204 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_205 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_205 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_206 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hce == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_206 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_207 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_207 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_208 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_208 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_209 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_209 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_210 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_210 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_211 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_211 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_212 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_212 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_213 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_213 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_214 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_214 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_215 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_215 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_216 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_216 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_217 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_217 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_218 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hda == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_218 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_219 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_219 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_220 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_220 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_221 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_221 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_222 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hde == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_222 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_223 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_223 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_224 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_224 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_225 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_225 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_226 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_226 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_227 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_227 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_228 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_228 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_229 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_229 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_230 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_230 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_231 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_231 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_232 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_232 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_233 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_233 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_234 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hea == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_234 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_235 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'heb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_235 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_236 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hec == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_236 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_237 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hed == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_237 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_238 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hee == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_238 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_239 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hef == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_239 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_240 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_240 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_241 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_241 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_242 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_242 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_243 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_243 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_244 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_244 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_245 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_245 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_246 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_246 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_247 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_247 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_248 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_248 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_249 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_249 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_250 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfa == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_250 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_251 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_251 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_252 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_252 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_253 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_253 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_254 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfe == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_254 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_255 <= 2'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hff == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_255 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (8'hff == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_255; // @[RAMWrapper.scala 43:22]
    end else if (8'hfe == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_254; // @[RAMWrapper.scala 43:22]
    end else if (8'hfd == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_253; // @[RAMWrapper.scala 43:22]
    end else if (8'hfc == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_252; // @[RAMWrapper.scala 43:22]
    end else begin
      io_douta_REG <= _GEN_251;
    end
    if (8'hff == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_255; // @[RAMWrapper.scala 44:22]
    end else if (8'hfe == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_254; // @[RAMWrapper.scala 44:22]
    end else if (8'hfd == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_253; // @[RAMWrapper.scala 44:22]
    end else if (8'hfc == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_252; // @[RAMWrapper.scala 44:22]
    end else begin
      io_doutb_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  mem_128 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  mem_129 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  mem_130 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  mem_131 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  mem_132 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  mem_133 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  mem_134 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  mem_135 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  mem_136 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  mem_137 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  mem_138 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  mem_139 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  mem_140 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  mem_141 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  mem_142 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  mem_143 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  mem_144 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  mem_145 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  mem_146 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  mem_147 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  mem_148 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  mem_149 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  mem_150 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  mem_151 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  mem_152 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  mem_153 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  mem_154 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  mem_155 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  mem_156 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  mem_157 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  mem_158 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  mem_159 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  mem_160 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  mem_161 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  mem_162 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  mem_163 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  mem_164 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  mem_165 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  mem_166 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  mem_167 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  mem_168 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  mem_169 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  mem_170 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  mem_171 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  mem_172 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  mem_173 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  mem_174 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  mem_175 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  mem_176 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  mem_177 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  mem_178 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  mem_179 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  mem_180 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  mem_181 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  mem_182 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  mem_183 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  mem_184 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  mem_185 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  mem_186 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  mem_187 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  mem_188 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  mem_189 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  mem_190 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  mem_191 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  mem_192 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  mem_193 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  mem_194 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  mem_195 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  mem_196 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  mem_197 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  mem_198 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  mem_199 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  mem_200 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  mem_201 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  mem_202 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  mem_203 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  mem_204 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  mem_205 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  mem_206 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  mem_207 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  mem_208 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  mem_209 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  mem_210 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  mem_211 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  mem_212 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  mem_213 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  mem_214 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  mem_215 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  mem_216 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  mem_217 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  mem_218 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  mem_219 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  mem_220 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  mem_221 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  mem_222 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  mem_223 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  mem_224 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  mem_225 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  mem_226 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  mem_227 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  mem_228 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  mem_229 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  mem_230 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  mem_231 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  mem_232 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  mem_233 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  mem_234 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  mem_235 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  mem_236 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  mem_237 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  mem_238 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  mem_239 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  mem_240 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  mem_241 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  mem_242 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  mem_243 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  mem_244 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  mem_245 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  mem_246 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  mem_247 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  mem_248 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  mem_249 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  mem_250 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  mem_251 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  mem_252 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  mem_253 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  mem_254 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  mem_255 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  io_douta_REG = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  io_doutb_REG = _RAND_257[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM(
  input        clock,
  input        reset,
  input        io_wea,
  input  [7:0] io_addra,
  input  [7:0] io_addrb,
  input  [1:0] io_dina,
  output [1:0] io_douta,
  output [1:0] io_doutb
);
  wire  sim_dual_port_bram_clock; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_reset; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_io_wea; // @[RAMWrapper.scala 30:36]
  wire [7:0] sim_dual_port_bram_io_addra; // @[RAMWrapper.scala 30:36]
  wire [7:0] sim_dual_port_bram_io_addrb; // @[RAMWrapper.scala 30:36]
  wire [1:0] sim_dual_port_bram_io_dina; // @[RAMWrapper.scala 30:36]
  wire [1:0] sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 30:36]
  wire [1:0] sim_dual_port_bram_io_doutb; // @[RAMWrapper.scala 30:36]
  SimDualPortBRAM sim_dual_port_bram ( // @[RAMWrapper.scala 30:36]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_wea(sim_dual_port_bram_io_wea),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dina(sim_dual_port_bram_io_dina),
    .io_douta(sim_dual_port_bram_io_douta),
    .io_doutb(sim_dual_port_bram_io_doutb)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 31:27]
  assign io_doutb = sim_dual_port_bram_io_doutb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_wea = io_wea; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_dina = io_dina; // @[RAMWrapper.scala 31:27]
endmodule
module SimDualPortBRAM_1(
  input         clock,
  input         reset,
  input         io_wea,
  input  [7:0]  io_addra,
  input  [7:0]  io_addrb,
  input  [61:0] io_dina,
  output [61:0] io_douta,
  output [61:0] io_doutb
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [63:0] _RAND_257;
`endif // RANDOMIZE_REG_INIT
  reg [61:0] mem_0; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_1; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_2; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_3; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_4; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_5; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_6; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_7; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_8; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_9; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_10; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_11; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_12; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_13; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_14; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_15; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_16; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_17; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_18; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_19; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_20; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_21; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_22; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_23; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_24; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_25; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_26; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_27; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_28; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_29; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_30; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_31; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_32; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_33; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_34; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_35; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_36; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_37; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_38; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_39; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_40; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_41; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_42; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_43; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_44; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_45; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_46; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_47; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_48; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_49; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_50; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_51; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_52; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_53; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_54; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_55; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_56; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_57; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_58; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_59; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_60; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_61; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_62; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_63; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_64; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_65; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_66; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_67; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_68; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_69; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_70; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_71; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_72; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_73; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_74; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_75; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_76; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_77; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_78; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_79; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_80; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_81; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_82; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_83; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_84; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_85; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_86; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_87; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_88; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_89; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_90; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_91; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_92; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_93; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_94; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_95; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_96; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_97; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_98; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_99; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_100; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_101; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_102; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_103; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_104; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_105; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_106; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_107; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_108; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_109; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_110; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_111; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_112; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_113; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_114; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_115; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_116; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_117; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_118; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_119; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_120; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_121; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_122; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_123; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_124; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_125; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_126; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_127; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_128; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_129; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_130; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_131; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_132; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_133; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_134; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_135; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_136; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_137; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_138; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_139; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_140; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_141; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_142; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_143; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_144; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_145; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_146; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_147; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_148; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_149; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_150; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_151; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_152; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_153; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_154; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_155; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_156; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_157; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_158; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_159; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_160; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_161; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_162; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_163; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_164; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_165; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_166; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_167; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_168; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_169; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_170; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_171; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_172; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_173; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_174; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_175; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_176; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_177; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_178; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_179; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_180; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_181; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_182; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_183; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_184; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_185; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_186; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_187; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_188; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_189; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_190; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_191; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_192; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_193; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_194; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_195; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_196; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_197; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_198; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_199; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_200; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_201; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_202; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_203; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_204; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_205; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_206; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_207; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_208; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_209; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_210; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_211; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_212; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_213; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_214; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_215; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_216; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_217; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_218; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_219; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_220; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_221; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_222; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_223; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_224; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_225; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_226; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_227; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_228; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_229; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_230; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_231; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_232; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_233; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_234; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_235; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_236; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_237; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_238; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_239; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_240; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_241; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_242; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_243; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_244; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_245; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_246; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_247; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_248; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_249; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_250; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_251; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_252; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_253; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_254; // @[RAMWrapper.scala 41:20]
  reg [61:0] mem_255; // @[RAMWrapper.scala 41:20]
  reg [61:0] io_douta_REG; // @[RAMWrapper.scala 43:22]
  wire [61:0] _GEN_1 = 8'h1 == io_addra ? mem_1 : mem_0; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_2 = 8'h2 == io_addra ? mem_2 : _GEN_1; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_3 = 8'h3 == io_addra ? mem_3 : _GEN_2; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_4 = 8'h4 == io_addra ? mem_4 : _GEN_3; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_5 = 8'h5 == io_addra ? mem_5 : _GEN_4; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_6 = 8'h6 == io_addra ? mem_6 : _GEN_5; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_7 = 8'h7 == io_addra ? mem_7 : _GEN_6; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_8 = 8'h8 == io_addra ? mem_8 : _GEN_7; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_9 = 8'h9 == io_addra ? mem_9 : _GEN_8; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_10 = 8'ha == io_addra ? mem_10 : _GEN_9; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_11 = 8'hb == io_addra ? mem_11 : _GEN_10; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_12 = 8'hc == io_addra ? mem_12 : _GEN_11; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_13 = 8'hd == io_addra ? mem_13 : _GEN_12; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_14 = 8'he == io_addra ? mem_14 : _GEN_13; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_15 = 8'hf == io_addra ? mem_15 : _GEN_14; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_16 = 8'h10 == io_addra ? mem_16 : _GEN_15; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_17 = 8'h11 == io_addra ? mem_17 : _GEN_16; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_18 = 8'h12 == io_addra ? mem_18 : _GEN_17; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_19 = 8'h13 == io_addra ? mem_19 : _GEN_18; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_20 = 8'h14 == io_addra ? mem_20 : _GEN_19; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_21 = 8'h15 == io_addra ? mem_21 : _GEN_20; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_22 = 8'h16 == io_addra ? mem_22 : _GEN_21; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_23 = 8'h17 == io_addra ? mem_23 : _GEN_22; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_24 = 8'h18 == io_addra ? mem_24 : _GEN_23; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_25 = 8'h19 == io_addra ? mem_25 : _GEN_24; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_26 = 8'h1a == io_addra ? mem_26 : _GEN_25; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_27 = 8'h1b == io_addra ? mem_27 : _GEN_26; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_28 = 8'h1c == io_addra ? mem_28 : _GEN_27; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_29 = 8'h1d == io_addra ? mem_29 : _GEN_28; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_30 = 8'h1e == io_addra ? mem_30 : _GEN_29; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_31 = 8'h1f == io_addra ? mem_31 : _GEN_30; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_32 = 8'h20 == io_addra ? mem_32 : _GEN_31; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_33 = 8'h21 == io_addra ? mem_33 : _GEN_32; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_34 = 8'h22 == io_addra ? mem_34 : _GEN_33; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_35 = 8'h23 == io_addra ? mem_35 : _GEN_34; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_36 = 8'h24 == io_addra ? mem_36 : _GEN_35; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_37 = 8'h25 == io_addra ? mem_37 : _GEN_36; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_38 = 8'h26 == io_addra ? mem_38 : _GEN_37; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_39 = 8'h27 == io_addra ? mem_39 : _GEN_38; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_40 = 8'h28 == io_addra ? mem_40 : _GEN_39; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_41 = 8'h29 == io_addra ? mem_41 : _GEN_40; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_42 = 8'h2a == io_addra ? mem_42 : _GEN_41; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_43 = 8'h2b == io_addra ? mem_43 : _GEN_42; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_44 = 8'h2c == io_addra ? mem_44 : _GEN_43; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_45 = 8'h2d == io_addra ? mem_45 : _GEN_44; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_46 = 8'h2e == io_addra ? mem_46 : _GEN_45; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_47 = 8'h2f == io_addra ? mem_47 : _GEN_46; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_48 = 8'h30 == io_addra ? mem_48 : _GEN_47; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_49 = 8'h31 == io_addra ? mem_49 : _GEN_48; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_50 = 8'h32 == io_addra ? mem_50 : _GEN_49; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_51 = 8'h33 == io_addra ? mem_51 : _GEN_50; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_52 = 8'h34 == io_addra ? mem_52 : _GEN_51; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_53 = 8'h35 == io_addra ? mem_53 : _GEN_52; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_54 = 8'h36 == io_addra ? mem_54 : _GEN_53; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_55 = 8'h37 == io_addra ? mem_55 : _GEN_54; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_56 = 8'h38 == io_addra ? mem_56 : _GEN_55; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_57 = 8'h39 == io_addra ? mem_57 : _GEN_56; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_58 = 8'h3a == io_addra ? mem_58 : _GEN_57; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_59 = 8'h3b == io_addra ? mem_59 : _GEN_58; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_60 = 8'h3c == io_addra ? mem_60 : _GEN_59; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_61 = 8'h3d == io_addra ? mem_61 : _GEN_60; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_62 = 8'h3e == io_addra ? mem_62 : _GEN_61; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_63 = 8'h3f == io_addra ? mem_63 : _GEN_62; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_64 = 8'h40 == io_addra ? mem_64 : _GEN_63; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_65 = 8'h41 == io_addra ? mem_65 : _GEN_64; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_66 = 8'h42 == io_addra ? mem_66 : _GEN_65; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_67 = 8'h43 == io_addra ? mem_67 : _GEN_66; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_68 = 8'h44 == io_addra ? mem_68 : _GEN_67; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_69 = 8'h45 == io_addra ? mem_69 : _GEN_68; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_70 = 8'h46 == io_addra ? mem_70 : _GEN_69; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_71 = 8'h47 == io_addra ? mem_71 : _GEN_70; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_72 = 8'h48 == io_addra ? mem_72 : _GEN_71; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_73 = 8'h49 == io_addra ? mem_73 : _GEN_72; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_74 = 8'h4a == io_addra ? mem_74 : _GEN_73; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_75 = 8'h4b == io_addra ? mem_75 : _GEN_74; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_76 = 8'h4c == io_addra ? mem_76 : _GEN_75; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_77 = 8'h4d == io_addra ? mem_77 : _GEN_76; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_78 = 8'h4e == io_addra ? mem_78 : _GEN_77; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_79 = 8'h4f == io_addra ? mem_79 : _GEN_78; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_80 = 8'h50 == io_addra ? mem_80 : _GEN_79; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_81 = 8'h51 == io_addra ? mem_81 : _GEN_80; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_82 = 8'h52 == io_addra ? mem_82 : _GEN_81; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_83 = 8'h53 == io_addra ? mem_83 : _GEN_82; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_84 = 8'h54 == io_addra ? mem_84 : _GEN_83; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_85 = 8'h55 == io_addra ? mem_85 : _GEN_84; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_86 = 8'h56 == io_addra ? mem_86 : _GEN_85; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_87 = 8'h57 == io_addra ? mem_87 : _GEN_86; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_88 = 8'h58 == io_addra ? mem_88 : _GEN_87; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_89 = 8'h59 == io_addra ? mem_89 : _GEN_88; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_90 = 8'h5a == io_addra ? mem_90 : _GEN_89; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_91 = 8'h5b == io_addra ? mem_91 : _GEN_90; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_92 = 8'h5c == io_addra ? mem_92 : _GEN_91; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_93 = 8'h5d == io_addra ? mem_93 : _GEN_92; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_94 = 8'h5e == io_addra ? mem_94 : _GEN_93; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_95 = 8'h5f == io_addra ? mem_95 : _GEN_94; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_96 = 8'h60 == io_addra ? mem_96 : _GEN_95; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_97 = 8'h61 == io_addra ? mem_97 : _GEN_96; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_98 = 8'h62 == io_addra ? mem_98 : _GEN_97; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_99 = 8'h63 == io_addra ? mem_99 : _GEN_98; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_100 = 8'h64 == io_addra ? mem_100 : _GEN_99; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_101 = 8'h65 == io_addra ? mem_101 : _GEN_100; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_102 = 8'h66 == io_addra ? mem_102 : _GEN_101; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_103 = 8'h67 == io_addra ? mem_103 : _GEN_102; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_104 = 8'h68 == io_addra ? mem_104 : _GEN_103; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_105 = 8'h69 == io_addra ? mem_105 : _GEN_104; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_106 = 8'h6a == io_addra ? mem_106 : _GEN_105; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_107 = 8'h6b == io_addra ? mem_107 : _GEN_106; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_108 = 8'h6c == io_addra ? mem_108 : _GEN_107; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_109 = 8'h6d == io_addra ? mem_109 : _GEN_108; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_110 = 8'h6e == io_addra ? mem_110 : _GEN_109; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_111 = 8'h6f == io_addra ? mem_111 : _GEN_110; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_112 = 8'h70 == io_addra ? mem_112 : _GEN_111; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_113 = 8'h71 == io_addra ? mem_113 : _GEN_112; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_114 = 8'h72 == io_addra ? mem_114 : _GEN_113; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_115 = 8'h73 == io_addra ? mem_115 : _GEN_114; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_116 = 8'h74 == io_addra ? mem_116 : _GEN_115; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_117 = 8'h75 == io_addra ? mem_117 : _GEN_116; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_118 = 8'h76 == io_addra ? mem_118 : _GEN_117; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_119 = 8'h77 == io_addra ? mem_119 : _GEN_118; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_120 = 8'h78 == io_addra ? mem_120 : _GEN_119; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_121 = 8'h79 == io_addra ? mem_121 : _GEN_120; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_122 = 8'h7a == io_addra ? mem_122 : _GEN_121; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_123 = 8'h7b == io_addra ? mem_123 : _GEN_122; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_124 = 8'h7c == io_addra ? mem_124 : _GEN_123; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_125 = 8'h7d == io_addra ? mem_125 : _GEN_124; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_126 = 8'h7e == io_addra ? mem_126 : _GEN_125; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_127 = 8'h7f == io_addra ? mem_127 : _GEN_126; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_128 = 8'h80 == io_addra ? mem_128 : _GEN_127; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_129 = 8'h81 == io_addra ? mem_129 : _GEN_128; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_130 = 8'h82 == io_addra ? mem_130 : _GEN_129; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_131 = 8'h83 == io_addra ? mem_131 : _GEN_130; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_132 = 8'h84 == io_addra ? mem_132 : _GEN_131; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_133 = 8'h85 == io_addra ? mem_133 : _GEN_132; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_134 = 8'h86 == io_addra ? mem_134 : _GEN_133; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_135 = 8'h87 == io_addra ? mem_135 : _GEN_134; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_136 = 8'h88 == io_addra ? mem_136 : _GEN_135; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_137 = 8'h89 == io_addra ? mem_137 : _GEN_136; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_138 = 8'h8a == io_addra ? mem_138 : _GEN_137; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_139 = 8'h8b == io_addra ? mem_139 : _GEN_138; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_140 = 8'h8c == io_addra ? mem_140 : _GEN_139; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_141 = 8'h8d == io_addra ? mem_141 : _GEN_140; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_142 = 8'h8e == io_addra ? mem_142 : _GEN_141; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_143 = 8'h8f == io_addra ? mem_143 : _GEN_142; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_144 = 8'h90 == io_addra ? mem_144 : _GEN_143; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_145 = 8'h91 == io_addra ? mem_145 : _GEN_144; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_146 = 8'h92 == io_addra ? mem_146 : _GEN_145; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_147 = 8'h93 == io_addra ? mem_147 : _GEN_146; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_148 = 8'h94 == io_addra ? mem_148 : _GEN_147; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_149 = 8'h95 == io_addra ? mem_149 : _GEN_148; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_150 = 8'h96 == io_addra ? mem_150 : _GEN_149; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_151 = 8'h97 == io_addra ? mem_151 : _GEN_150; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_152 = 8'h98 == io_addra ? mem_152 : _GEN_151; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_153 = 8'h99 == io_addra ? mem_153 : _GEN_152; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_154 = 8'h9a == io_addra ? mem_154 : _GEN_153; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_155 = 8'h9b == io_addra ? mem_155 : _GEN_154; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_156 = 8'h9c == io_addra ? mem_156 : _GEN_155; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_157 = 8'h9d == io_addra ? mem_157 : _GEN_156; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_158 = 8'h9e == io_addra ? mem_158 : _GEN_157; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_159 = 8'h9f == io_addra ? mem_159 : _GEN_158; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_160 = 8'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_161 = 8'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_162 = 8'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_163 = 8'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_164 = 8'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_165 = 8'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_166 = 8'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_167 = 8'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_168 = 8'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_169 = 8'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_170 = 8'haa == io_addra ? mem_170 : _GEN_169; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_171 = 8'hab == io_addra ? mem_171 : _GEN_170; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_172 = 8'hac == io_addra ? mem_172 : _GEN_171; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_173 = 8'had == io_addra ? mem_173 : _GEN_172; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_174 = 8'hae == io_addra ? mem_174 : _GEN_173; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_175 = 8'haf == io_addra ? mem_175 : _GEN_174; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_176 = 8'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_177 = 8'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_178 = 8'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_179 = 8'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_180 = 8'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_181 = 8'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_182 = 8'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_183 = 8'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_184 = 8'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_185 = 8'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_186 = 8'hba == io_addra ? mem_186 : _GEN_185; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_187 = 8'hbb == io_addra ? mem_187 : _GEN_186; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_188 = 8'hbc == io_addra ? mem_188 : _GEN_187; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_189 = 8'hbd == io_addra ? mem_189 : _GEN_188; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_190 = 8'hbe == io_addra ? mem_190 : _GEN_189; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_191 = 8'hbf == io_addra ? mem_191 : _GEN_190; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_192 = 8'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_193 = 8'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_194 = 8'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_195 = 8'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_196 = 8'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_197 = 8'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_198 = 8'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_199 = 8'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_200 = 8'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_201 = 8'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_202 = 8'hca == io_addra ? mem_202 : _GEN_201; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_203 = 8'hcb == io_addra ? mem_203 : _GEN_202; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_204 = 8'hcc == io_addra ? mem_204 : _GEN_203; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_205 = 8'hcd == io_addra ? mem_205 : _GEN_204; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_206 = 8'hce == io_addra ? mem_206 : _GEN_205; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_207 = 8'hcf == io_addra ? mem_207 : _GEN_206; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_208 = 8'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_209 = 8'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_210 = 8'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_211 = 8'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_212 = 8'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_213 = 8'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_214 = 8'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_215 = 8'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_216 = 8'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_217 = 8'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_218 = 8'hda == io_addra ? mem_218 : _GEN_217; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_219 = 8'hdb == io_addra ? mem_219 : _GEN_218; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_220 = 8'hdc == io_addra ? mem_220 : _GEN_219; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_221 = 8'hdd == io_addra ? mem_221 : _GEN_220; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_222 = 8'hde == io_addra ? mem_222 : _GEN_221; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_223 = 8'hdf == io_addra ? mem_223 : _GEN_222; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_224 = 8'he0 == io_addra ? mem_224 : _GEN_223; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_225 = 8'he1 == io_addra ? mem_225 : _GEN_224; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_226 = 8'he2 == io_addra ? mem_226 : _GEN_225; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_227 = 8'he3 == io_addra ? mem_227 : _GEN_226; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_228 = 8'he4 == io_addra ? mem_228 : _GEN_227; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_229 = 8'he5 == io_addra ? mem_229 : _GEN_228; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_230 = 8'he6 == io_addra ? mem_230 : _GEN_229; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_231 = 8'he7 == io_addra ? mem_231 : _GEN_230; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_232 = 8'he8 == io_addra ? mem_232 : _GEN_231; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_233 = 8'he9 == io_addra ? mem_233 : _GEN_232; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_234 = 8'hea == io_addra ? mem_234 : _GEN_233; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_235 = 8'heb == io_addra ? mem_235 : _GEN_234; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_236 = 8'hec == io_addra ? mem_236 : _GEN_235; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_237 = 8'hed == io_addra ? mem_237 : _GEN_236; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_238 = 8'hee == io_addra ? mem_238 : _GEN_237; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_239 = 8'hef == io_addra ? mem_239 : _GEN_238; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_240 = 8'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_241 = 8'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_242 = 8'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_243 = 8'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_244 = 8'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_245 = 8'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_246 = 8'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_247 = 8'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_248 = 8'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_249 = 8'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_250 = 8'hfa == io_addra ? mem_250 : _GEN_249; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [61:0] _GEN_251 = 8'hfb == io_addra ? mem_251 : _GEN_250; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  reg [61:0] io_doutb_REG; // @[RAMWrapper.scala 44:22]
  wire [61:0] _GEN_257 = 8'h1 == io_addrb ? mem_1 : mem_0; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_258 = 8'h2 == io_addrb ? mem_2 : _GEN_257; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_259 = 8'h3 == io_addrb ? mem_3 : _GEN_258; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_260 = 8'h4 == io_addrb ? mem_4 : _GEN_259; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_261 = 8'h5 == io_addrb ? mem_5 : _GEN_260; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_262 = 8'h6 == io_addrb ? mem_6 : _GEN_261; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_263 = 8'h7 == io_addrb ? mem_7 : _GEN_262; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_264 = 8'h8 == io_addrb ? mem_8 : _GEN_263; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_265 = 8'h9 == io_addrb ? mem_9 : _GEN_264; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_266 = 8'ha == io_addrb ? mem_10 : _GEN_265; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_267 = 8'hb == io_addrb ? mem_11 : _GEN_266; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_268 = 8'hc == io_addrb ? mem_12 : _GEN_267; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_269 = 8'hd == io_addrb ? mem_13 : _GEN_268; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_270 = 8'he == io_addrb ? mem_14 : _GEN_269; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_271 = 8'hf == io_addrb ? mem_15 : _GEN_270; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_272 = 8'h10 == io_addrb ? mem_16 : _GEN_271; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_273 = 8'h11 == io_addrb ? mem_17 : _GEN_272; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_274 = 8'h12 == io_addrb ? mem_18 : _GEN_273; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_275 = 8'h13 == io_addrb ? mem_19 : _GEN_274; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_276 = 8'h14 == io_addrb ? mem_20 : _GEN_275; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_277 = 8'h15 == io_addrb ? mem_21 : _GEN_276; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_278 = 8'h16 == io_addrb ? mem_22 : _GEN_277; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_279 = 8'h17 == io_addrb ? mem_23 : _GEN_278; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_280 = 8'h18 == io_addrb ? mem_24 : _GEN_279; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_281 = 8'h19 == io_addrb ? mem_25 : _GEN_280; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_282 = 8'h1a == io_addrb ? mem_26 : _GEN_281; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_283 = 8'h1b == io_addrb ? mem_27 : _GEN_282; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_284 = 8'h1c == io_addrb ? mem_28 : _GEN_283; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_285 = 8'h1d == io_addrb ? mem_29 : _GEN_284; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_286 = 8'h1e == io_addrb ? mem_30 : _GEN_285; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_287 = 8'h1f == io_addrb ? mem_31 : _GEN_286; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_288 = 8'h20 == io_addrb ? mem_32 : _GEN_287; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_289 = 8'h21 == io_addrb ? mem_33 : _GEN_288; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_290 = 8'h22 == io_addrb ? mem_34 : _GEN_289; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_291 = 8'h23 == io_addrb ? mem_35 : _GEN_290; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_292 = 8'h24 == io_addrb ? mem_36 : _GEN_291; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_293 = 8'h25 == io_addrb ? mem_37 : _GEN_292; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_294 = 8'h26 == io_addrb ? mem_38 : _GEN_293; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_295 = 8'h27 == io_addrb ? mem_39 : _GEN_294; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_296 = 8'h28 == io_addrb ? mem_40 : _GEN_295; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_297 = 8'h29 == io_addrb ? mem_41 : _GEN_296; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_298 = 8'h2a == io_addrb ? mem_42 : _GEN_297; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_299 = 8'h2b == io_addrb ? mem_43 : _GEN_298; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_300 = 8'h2c == io_addrb ? mem_44 : _GEN_299; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_301 = 8'h2d == io_addrb ? mem_45 : _GEN_300; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_302 = 8'h2e == io_addrb ? mem_46 : _GEN_301; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_303 = 8'h2f == io_addrb ? mem_47 : _GEN_302; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_304 = 8'h30 == io_addrb ? mem_48 : _GEN_303; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_305 = 8'h31 == io_addrb ? mem_49 : _GEN_304; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_306 = 8'h32 == io_addrb ? mem_50 : _GEN_305; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_307 = 8'h33 == io_addrb ? mem_51 : _GEN_306; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_308 = 8'h34 == io_addrb ? mem_52 : _GEN_307; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_309 = 8'h35 == io_addrb ? mem_53 : _GEN_308; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_310 = 8'h36 == io_addrb ? mem_54 : _GEN_309; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_311 = 8'h37 == io_addrb ? mem_55 : _GEN_310; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_312 = 8'h38 == io_addrb ? mem_56 : _GEN_311; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_313 = 8'h39 == io_addrb ? mem_57 : _GEN_312; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_314 = 8'h3a == io_addrb ? mem_58 : _GEN_313; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_315 = 8'h3b == io_addrb ? mem_59 : _GEN_314; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_316 = 8'h3c == io_addrb ? mem_60 : _GEN_315; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_317 = 8'h3d == io_addrb ? mem_61 : _GEN_316; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_318 = 8'h3e == io_addrb ? mem_62 : _GEN_317; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_319 = 8'h3f == io_addrb ? mem_63 : _GEN_318; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_320 = 8'h40 == io_addrb ? mem_64 : _GEN_319; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_321 = 8'h41 == io_addrb ? mem_65 : _GEN_320; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_322 = 8'h42 == io_addrb ? mem_66 : _GEN_321; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_323 = 8'h43 == io_addrb ? mem_67 : _GEN_322; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_324 = 8'h44 == io_addrb ? mem_68 : _GEN_323; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_325 = 8'h45 == io_addrb ? mem_69 : _GEN_324; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_326 = 8'h46 == io_addrb ? mem_70 : _GEN_325; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_327 = 8'h47 == io_addrb ? mem_71 : _GEN_326; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_328 = 8'h48 == io_addrb ? mem_72 : _GEN_327; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_329 = 8'h49 == io_addrb ? mem_73 : _GEN_328; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_330 = 8'h4a == io_addrb ? mem_74 : _GEN_329; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_331 = 8'h4b == io_addrb ? mem_75 : _GEN_330; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_332 = 8'h4c == io_addrb ? mem_76 : _GEN_331; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_333 = 8'h4d == io_addrb ? mem_77 : _GEN_332; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_334 = 8'h4e == io_addrb ? mem_78 : _GEN_333; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_335 = 8'h4f == io_addrb ? mem_79 : _GEN_334; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_336 = 8'h50 == io_addrb ? mem_80 : _GEN_335; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_337 = 8'h51 == io_addrb ? mem_81 : _GEN_336; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_338 = 8'h52 == io_addrb ? mem_82 : _GEN_337; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_339 = 8'h53 == io_addrb ? mem_83 : _GEN_338; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_340 = 8'h54 == io_addrb ? mem_84 : _GEN_339; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_341 = 8'h55 == io_addrb ? mem_85 : _GEN_340; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_342 = 8'h56 == io_addrb ? mem_86 : _GEN_341; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_343 = 8'h57 == io_addrb ? mem_87 : _GEN_342; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_344 = 8'h58 == io_addrb ? mem_88 : _GEN_343; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_345 = 8'h59 == io_addrb ? mem_89 : _GEN_344; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_346 = 8'h5a == io_addrb ? mem_90 : _GEN_345; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_347 = 8'h5b == io_addrb ? mem_91 : _GEN_346; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_348 = 8'h5c == io_addrb ? mem_92 : _GEN_347; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_349 = 8'h5d == io_addrb ? mem_93 : _GEN_348; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_350 = 8'h5e == io_addrb ? mem_94 : _GEN_349; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_351 = 8'h5f == io_addrb ? mem_95 : _GEN_350; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_352 = 8'h60 == io_addrb ? mem_96 : _GEN_351; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_353 = 8'h61 == io_addrb ? mem_97 : _GEN_352; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_354 = 8'h62 == io_addrb ? mem_98 : _GEN_353; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_355 = 8'h63 == io_addrb ? mem_99 : _GEN_354; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_356 = 8'h64 == io_addrb ? mem_100 : _GEN_355; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_357 = 8'h65 == io_addrb ? mem_101 : _GEN_356; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_358 = 8'h66 == io_addrb ? mem_102 : _GEN_357; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_359 = 8'h67 == io_addrb ? mem_103 : _GEN_358; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_360 = 8'h68 == io_addrb ? mem_104 : _GEN_359; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_361 = 8'h69 == io_addrb ? mem_105 : _GEN_360; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_362 = 8'h6a == io_addrb ? mem_106 : _GEN_361; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_363 = 8'h6b == io_addrb ? mem_107 : _GEN_362; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_364 = 8'h6c == io_addrb ? mem_108 : _GEN_363; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_365 = 8'h6d == io_addrb ? mem_109 : _GEN_364; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_366 = 8'h6e == io_addrb ? mem_110 : _GEN_365; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_367 = 8'h6f == io_addrb ? mem_111 : _GEN_366; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_368 = 8'h70 == io_addrb ? mem_112 : _GEN_367; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_369 = 8'h71 == io_addrb ? mem_113 : _GEN_368; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_370 = 8'h72 == io_addrb ? mem_114 : _GEN_369; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_371 = 8'h73 == io_addrb ? mem_115 : _GEN_370; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_372 = 8'h74 == io_addrb ? mem_116 : _GEN_371; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_373 = 8'h75 == io_addrb ? mem_117 : _GEN_372; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_374 = 8'h76 == io_addrb ? mem_118 : _GEN_373; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_375 = 8'h77 == io_addrb ? mem_119 : _GEN_374; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_376 = 8'h78 == io_addrb ? mem_120 : _GEN_375; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_377 = 8'h79 == io_addrb ? mem_121 : _GEN_376; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_378 = 8'h7a == io_addrb ? mem_122 : _GEN_377; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_379 = 8'h7b == io_addrb ? mem_123 : _GEN_378; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_380 = 8'h7c == io_addrb ? mem_124 : _GEN_379; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_381 = 8'h7d == io_addrb ? mem_125 : _GEN_380; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_382 = 8'h7e == io_addrb ? mem_126 : _GEN_381; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_383 = 8'h7f == io_addrb ? mem_127 : _GEN_382; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_384 = 8'h80 == io_addrb ? mem_128 : _GEN_383; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_385 = 8'h81 == io_addrb ? mem_129 : _GEN_384; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_386 = 8'h82 == io_addrb ? mem_130 : _GEN_385; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_387 = 8'h83 == io_addrb ? mem_131 : _GEN_386; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_388 = 8'h84 == io_addrb ? mem_132 : _GEN_387; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_389 = 8'h85 == io_addrb ? mem_133 : _GEN_388; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_390 = 8'h86 == io_addrb ? mem_134 : _GEN_389; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_391 = 8'h87 == io_addrb ? mem_135 : _GEN_390; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_392 = 8'h88 == io_addrb ? mem_136 : _GEN_391; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_393 = 8'h89 == io_addrb ? mem_137 : _GEN_392; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_394 = 8'h8a == io_addrb ? mem_138 : _GEN_393; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_395 = 8'h8b == io_addrb ? mem_139 : _GEN_394; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_396 = 8'h8c == io_addrb ? mem_140 : _GEN_395; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_397 = 8'h8d == io_addrb ? mem_141 : _GEN_396; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_398 = 8'h8e == io_addrb ? mem_142 : _GEN_397; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_399 = 8'h8f == io_addrb ? mem_143 : _GEN_398; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_400 = 8'h90 == io_addrb ? mem_144 : _GEN_399; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_401 = 8'h91 == io_addrb ? mem_145 : _GEN_400; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_402 = 8'h92 == io_addrb ? mem_146 : _GEN_401; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_403 = 8'h93 == io_addrb ? mem_147 : _GEN_402; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_404 = 8'h94 == io_addrb ? mem_148 : _GEN_403; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_405 = 8'h95 == io_addrb ? mem_149 : _GEN_404; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_406 = 8'h96 == io_addrb ? mem_150 : _GEN_405; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_407 = 8'h97 == io_addrb ? mem_151 : _GEN_406; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_408 = 8'h98 == io_addrb ? mem_152 : _GEN_407; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_409 = 8'h99 == io_addrb ? mem_153 : _GEN_408; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_410 = 8'h9a == io_addrb ? mem_154 : _GEN_409; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_411 = 8'h9b == io_addrb ? mem_155 : _GEN_410; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_412 = 8'h9c == io_addrb ? mem_156 : _GEN_411; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_413 = 8'h9d == io_addrb ? mem_157 : _GEN_412; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_414 = 8'h9e == io_addrb ? mem_158 : _GEN_413; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_415 = 8'h9f == io_addrb ? mem_159 : _GEN_414; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_416 = 8'ha0 == io_addrb ? mem_160 : _GEN_415; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_417 = 8'ha1 == io_addrb ? mem_161 : _GEN_416; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_418 = 8'ha2 == io_addrb ? mem_162 : _GEN_417; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_419 = 8'ha3 == io_addrb ? mem_163 : _GEN_418; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_420 = 8'ha4 == io_addrb ? mem_164 : _GEN_419; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_421 = 8'ha5 == io_addrb ? mem_165 : _GEN_420; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_422 = 8'ha6 == io_addrb ? mem_166 : _GEN_421; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_423 = 8'ha7 == io_addrb ? mem_167 : _GEN_422; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_424 = 8'ha8 == io_addrb ? mem_168 : _GEN_423; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_425 = 8'ha9 == io_addrb ? mem_169 : _GEN_424; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_426 = 8'haa == io_addrb ? mem_170 : _GEN_425; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_427 = 8'hab == io_addrb ? mem_171 : _GEN_426; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_428 = 8'hac == io_addrb ? mem_172 : _GEN_427; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_429 = 8'had == io_addrb ? mem_173 : _GEN_428; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_430 = 8'hae == io_addrb ? mem_174 : _GEN_429; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_431 = 8'haf == io_addrb ? mem_175 : _GEN_430; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_432 = 8'hb0 == io_addrb ? mem_176 : _GEN_431; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_433 = 8'hb1 == io_addrb ? mem_177 : _GEN_432; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_434 = 8'hb2 == io_addrb ? mem_178 : _GEN_433; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_435 = 8'hb3 == io_addrb ? mem_179 : _GEN_434; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_436 = 8'hb4 == io_addrb ? mem_180 : _GEN_435; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_437 = 8'hb5 == io_addrb ? mem_181 : _GEN_436; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_438 = 8'hb6 == io_addrb ? mem_182 : _GEN_437; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_439 = 8'hb7 == io_addrb ? mem_183 : _GEN_438; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_440 = 8'hb8 == io_addrb ? mem_184 : _GEN_439; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_441 = 8'hb9 == io_addrb ? mem_185 : _GEN_440; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_442 = 8'hba == io_addrb ? mem_186 : _GEN_441; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_443 = 8'hbb == io_addrb ? mem_187 : _GEN_442; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_444 = 8'hbc == io_addrb ? mem_188 : _GEN_443; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_445 = 8'hbd == io_addrb ? mem_189 : _GEN_444; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_446 = 8'hbe == io_addrb ? mem_190 : _GEN_445; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_447 = 8'hbf == io_addrb ? mem_191 : _GEN_446; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_448 = 8'hc0 == io_addrb ? mem_192 : _GEN_447; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_449 = 8'hc1 == io_addrb ? mem_193 : _GEN_448; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_450 = 8'hc2 == io_addrb ? mem_194 : _GEN_449; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_451 = 8'hc3 == io_addrb ? mem_195 : _GEN_450; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_452 = 8'hc4 == io_addrb ? mem_196 : _GEN_451; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_453 = 8'hc5 == io_addrb ? mem_197 : _GEN_452; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_454 = 8'hc6 == io_addrb ? mem_198 : _GEN_453; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_455 = 8'hc7 == io_addrb ? mem_199 : _GEN_454; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_456 = 8'hc8 == io_addrb ? mem_200 : _GEN_455; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_457 = 8'hc9 == io_addrb ? mem_201 : _GEN_456; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_458 = 8'hca == io_addrb ? mem_202 : _GEN_457; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_459 = 8'hcb == io_addrb ? mem_203 : _GEN_458; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_460 = 8'hcc == io_addrb ? mem_204 : _GEN_459; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_461 = 8'hcd == io_addrb ? mem_205 : _GEN_460; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_462 = 8'hce == io_addrb ? mem_206 : _GEN_461; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_463 = 8'hcf == io_addrb ? mem_207 : _GEN_462; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_464 = 8'hd0 == io_addrb ? mem_208 : _GEN_463; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_465 = 8'hd1 == io_addrb ? mem_209 : _GEN_464; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_466 = 8'hd2 == io_addrb ? mem_210 : _GEN_465; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_467 = 8'hd3 == io_addrb ? mem_211 : _GEN_466; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_468 = 8'hd4 == io_addrb ? mem_212 : _GEN_467; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_469 = 8'hd5 == io_addrb ? mem_213 : _GEN_468; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_470 = 8'hd6 == io_addrb ? mem_214 : _GEN_469; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_471 = 8'hd7 == io_addrb ? mem_215 : _GEN_470; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_472 = 8'hd8 == io_addrb ? mem_216 : _GEN_471; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_473 = 8'hd9 == io_addrb ? mem_217 : _GEN_472; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_474 = 8'hda == io_addrb ? mem_218 : _GEN_473; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_475 = 8'hdb == io_addrb ? mem_219 : _GEN_474; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_476 = 8'hdc == io_addrb ? mem_220 : _GEN_475; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_477 = 8'hdd == io_addrb ? mem_221 : _GEN_476; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_478 = 8'hde == io_addrb ? mem_222 : _GEN_477; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_479 = 8'hdf == io_addrb ? mem_223 : _GEN_478; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_480 = 8'he0 == io_addrb ? mem_224 : _GEN_479; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_481 = 8'he1 == io_addrb ? mem_225 : _GEN_480; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_482 = 8'he2 == io_addrb ? mem_226 : _GEN_481; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_483 = 8'he3 == io_addrb ? mem_227 : _GEN_482; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_484 = 8'he4 == io_addrb ? mem_228 : _GEN_483; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_485 = 8'he5 == io_addrb ? mem_229 : _GEN_484; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_486 = 8'he6 == io_addrb ? mem_230 : _GEN_485; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_487 = 8'he7 == io_addrb ? mem_231 : _GEN_486; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_488 = 8'he8 == io_addrb ? mem_232 : _GEN_487; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_489 = 8'he9 == io_addrb ? mem_233 : _GEN_488; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_490 = 8'hea == io_addrb ? mem_234 : _GEN_489; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_491 = 8'heb == io_addrb ? mem_235 : _GEN_490; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_492 = 8'hec == io_addrb ? mem_236 : _GEN_491; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_493 = 8'hed == io_addrb ? mem_237 : _GEN_492; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_494 = 8'hee == io_addrb ? mem_238 : _GEN_493; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_495 = 8'hef == io_addrb ? mem_239 : _GEN_494; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_496 = 8'hf0 == io_addrb ? mem_240 : _GEN_495; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_497 = 8'hf1 == io_addrb ? mem_241 : _GEN_496; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_498 = 8'hf2 == io_addrb ? mem_242 : _GEN_497; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_499 = 8'hf3 == io_addrb ? mem_243 : _GEN_498; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_500 = 8'hf4 == io_addrb ? mem_244 : _GEN_499; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_501 = 8'hf5 == io_addrb ? mem_245 : _GEN_500; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_502 = 8'hf6 == io_addrb ? mem_246 : _GEN_501; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_503 = 8'hf7 == io_addrb ? mem_247 : _GEN_502; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_504 = 8'hf8 == io_addrb ? mem_248 : _GEN_503; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_505 = 8'hf9 == io_addrb ? mem_249 : _GEN_504; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_506 = 8'hfa == io_addrb ? mem_250 : _GEN_505; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  wire [61:0] _GEN_507 = 8'hfb == io_addrb ? mem_251 : _GEN_506; // @[RAMWrapper.scala 44:22 RAMWrapper.scala 44:22]
  assign io_douta = io_douta_REG; // @[RAMWrapper.scala 43:12]
  assign io_doutb = io_doutb_REG; // @[RAMWrapper.scala 44:12]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_0 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_0 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_1 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_1 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_2 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_2 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_3 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_3 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_4 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_4 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_5 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_5 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_6 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_6 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_7 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_7 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_8 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_8 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_9 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_9 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_10 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_10 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_11 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_11 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_12 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_12 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_13 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_13 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_14 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_14 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_15 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_15 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_16 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h10 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_16 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_17 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h11 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_17 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_18 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h12 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_18 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_19 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h13 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_19 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_20 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h14 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_20 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_21 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h15 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_21 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_22 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h16 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_22 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_23 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h17 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_23 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_24 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h18 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_24 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_25 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h19 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_25 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_26 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_26 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_27 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_27 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_28 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_28 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_29 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_29 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_30 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_30 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_31 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h1f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_31 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_32 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h20 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_32 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_33 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h21 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_33 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_34 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h22 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_34 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_35 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h23 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_35 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_36 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h24 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_36 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_37 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h25 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_37 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_38 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h26 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_38 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_39 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h27 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_39 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_40 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h28 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_40 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_41 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h29 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_41 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_42 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_42 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_43 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_43 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_44 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_44 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_45 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_45 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_46 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_46 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_47 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h2f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_47 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_48 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h30 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_48 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_49 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h31 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_49 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_50 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h32 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_50 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_51 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h33 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_51 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_52 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h34 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_52 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_53 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h35 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_53 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_54 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h36 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_54 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_55 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h37 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_55 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_56 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h38 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_56 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_57 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h39 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_57 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_58 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_58 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_59 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_59 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_60 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_60 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_61 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_61 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_62 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_62 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_63 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h3f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_63 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_64 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h40 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_64 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_65 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h41 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_65 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_66 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h42 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_66 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_67 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h43 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_67 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_68 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h44 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_68 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_69 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h45 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_69 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_70 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h46 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_70 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_71 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h47 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_71 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_72 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h48 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_72 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_73 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h49 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_73 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_74 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_74 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_75 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_75 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_76 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_76 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_77 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_77 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_78 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_78 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_79 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h4f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_79 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_80 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h50 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_80 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_81 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h51 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_81 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_82 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h52 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_82 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_83 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h53 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_83 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_84 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h54 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_84 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_85 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h55 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_85 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_86 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h56 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_86 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_87 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h57 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_87 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_88 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h58 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_88 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_89 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h59 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_89 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_90 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_90 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_91 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_91 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_92 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_92 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_93 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_93 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_94 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_94 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_95 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h5f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_95 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_96 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h60 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_96 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_97 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h61 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_97 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_98 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h62 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_98 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_99 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h63 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_99 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_100 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h64 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_100 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_101 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h65 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_101 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_102 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h66 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_102 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_103 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h67 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_103 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_104 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h68 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_104 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_105 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h69 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_105 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_106 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_106 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_107 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_107 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_108 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_108 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_109 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_109 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_110 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_110 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_111 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h6f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_111 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_112 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h70 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_112 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_113 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h71 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_113 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_114 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h72 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_114 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_115 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h73 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_115 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_116 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h74 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_116 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_117 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h75 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_117 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_118 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h76 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_118 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_119 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h77 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_119 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_120 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h78 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_120 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_121 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h79 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_121 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_122 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_122 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_123 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_123 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_124 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_124 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_125 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_125 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_126 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_126 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_127 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h7f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_127 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_128 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h80 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_128 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_129 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h81 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_129 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_130 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h82 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_130 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_131 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h83 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_131 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_132 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h84 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_132 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_133 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h85 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_133 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_134 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h86 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_134 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_135 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h87 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_135 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_136 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h88 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_136 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_137 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h89 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_137 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_138 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_138 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_139 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_139 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_140 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_140 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_141 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_141 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_142 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_142 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_143 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h8f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_143 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_144 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h90 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_144 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_145 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h91 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_145 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_146 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h92 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_146 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_147 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h93 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_147 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_148 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h94 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_148 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_149 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h95 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_149 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_150 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h96 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_150 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_151 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h97 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_151 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_152 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h98 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_152 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_153 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h99 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_153 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_154 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9a == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_154 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_155 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9b == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_155 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_156 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9c == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_156 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_157 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9d == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_157 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_158 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9e == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_158 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_159 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'h9f == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_159 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_160 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_160 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_161 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_161 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_162 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_162 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_163 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_163 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_164 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_164 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_165 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_165 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_166 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_166 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_167 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_167 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_168 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_168 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_169 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'ha9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_169 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_170 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'haa == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_170 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_171 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hab == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_171 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_172 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hac == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_172 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_173 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'had == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_173 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_174 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hae == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_174 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_175 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'haf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_175 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_176 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_176 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_177 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_177 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_178 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_178 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_179 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_179 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_180 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_180 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_181 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_181 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_182 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_182 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_183 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_183 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_184 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_184 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_185 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hb9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_185 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_186 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hba == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_186 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_187 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_187 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_188 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_188 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_189 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_189 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_190 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbe == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_190 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_191 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hbf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_191 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_192 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_192 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_193 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_193 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_194 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_194 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_195 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_195 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_196 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_196 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_197 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_197 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_198 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_198 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_199 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_199 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_200 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_200 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_201 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hc9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_201 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_202 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hca == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_202 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_203 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_203 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_204 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_204 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_205 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_205 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_206 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hce == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_206 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_207 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hcf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_207 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_208 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_208 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_209 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_209 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_210 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_210 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_211 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_211 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_212 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_212 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_213 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_213 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_214 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_214 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_215 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_215 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_216 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_216 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_217 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hd9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_217 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_218 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hda == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_218 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_219 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_219 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_220 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_220 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_221 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_221 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_222 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hde == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_222 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_223 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hdf == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_223 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_224 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_224 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_225 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_225 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_226 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_226 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_227 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_227 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_228 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_228 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_229 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_229 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_230 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_230 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_231 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_231 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_232 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_232 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_233 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'he9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_233 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_234 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hea == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_234 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_235 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'heb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_235 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_236 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hec == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_236 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_237 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hed == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_237 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_238 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hee == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_238 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_239 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hef == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_239 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_240 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf0 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_240 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_241 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf1 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_241 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_242 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf2 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_242 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_243 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf3 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_243 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_244 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf4 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_244 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_245 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf5 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_245 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_246 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf6 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_246 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_247 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf7 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_247 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_248 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf8 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_248 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_249 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hf9 == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_249 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_250 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfa == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_250 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_251 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfb == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_251 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_252 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfc == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_252 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_253 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfd == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_253 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_254 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hfe == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_254 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_255 <= 62'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_wea) begin // @[RAMWrapper.scala 46:16]
      if (8'hff == io_addra) begin // @[RAMWrapper.scala 47:19]
        mem_255 <= io_dina; // @[RAMWrapper.scala 47:19]
      end
    end
    if (8'hff == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_255; // @[RAMWrapper.scala 43:22]
    end else if (8'hfe == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_254; // @[RAMWrapper.scala 43:22]
    end else if (8'hfd == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_253; // @[RAMWrapper.scala 43:22]
    end else if (8'hfc == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_252; // @[RAMWrapper.scala 43:22]
    end else begin
      io_douta_REG <= _GEN_251;
    end
    if (8'hff == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_255; // @[RAMWrapper.scala 44:22]
    end else if (8'hfe == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_254; // @[RAMWrapper.scala 44:22]
    end else if (8'hfd == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_253; // @[RAMWrapper.scala 44:22]
    end else if (8'hfc == io_addrb) begin // @[RAMWrapper.scala 44:22]
      io_doutb_REG <= mem_252; // @[RAMWrapper.scala 44:22]
    end else begin
      io_doutb_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mem_0 = _RAND_0[61:0];
  _RAND_1 = {2{`RANDOM}};
  mem_1 = _RAND_1[61:0];
  _RAND_2 = {2{`RANDOM}};
  mem_2 = _RAND_2[61:0];
  _RAND_3 = {2{`RANDOM}};
  mem_3 = _RAND_3[61:0];
  _RAND_4 = {2{`RANDOM}};
  mem_4 = _RAND_4[61:0];
  _RAND_5 = {2{`RANDOM}};
  mem_5 = _RAND_5[61:0];
  _RAND_6 = {2{`RANDOM}};
  mem_6 = _RAND_6[61:0];
  _RAND_7 = {2{`RANDOM}};
  mem_7 = _RAND_7[61:0];
  _RAND_8 = {2{`RANDOM}};
  mem_8 = _RAND_8[61:0];
  _RAND_9 = {2{`RANDOM}};
  mem_9 = _RAND_9[61:0];
  _RAND_10 = {2{`RANDOM}};
  mem_10 = _RAND_10[61:0];
  _RAND_11 = {2{`RANDOM}};
  mem_11 = _RAND_11[61:0];
  _RAND_12 = {2{`RANDOM}};
  mem_12 = _RAND_12[61:0];
  _RAND_13 = {2{`RANDOM}};
  mem_13 = _RAND_13[61:0];
  _RAND_14 = {2{`RANDOM}};
  mem_14 = _RAND_14[61:0];
  _RAND_15 = {2{`RANDOM}};
  mem_15 = _RAND_15[61:0];
  _RAND_16 = {2{`RANDOM}};
  mem_16 = _RAND_16[61:0];
  _RAND_17 = {2{`RANDOM}};
  mem_17 = _RAND_17[61:0];
  _RAND_18 = {2{`RANDOM}};
  mem_18 = _RAND_18[61:0];
  _RAND_19 = {2{`RANDOM}};
  mem_19 = _RAND_19[61:0];
  _RAND_20 = {2{`RANDOM}};
  mem_20 = _RAND_20[61:0];
  _RAND_21 = {2{`RANDOM}};
  mem_21 = _RAND_21[61:0];
  _RAND_22 = {2{`RANDOM}};
  mem_22 = _RAND_22[61:0];
  _RAND_23 = {2{`RANDOM}};
  mem_23 = _RAND_23[61:0];
  _RAND_24 = {2{`RANDOM}};
  mem_24 = _RAND_24[61:0];
  _RAND_25 = {2{`RANDOM}};
  mem_25 = _RAND_25[61:0];
  _RAND_26 = {2{`RANDOM}};
  mem_26 = _RAND_26[61:0];
  _RAND_27 = {2{`RANDOM}};
  mem_27 = _RAND_27[61:0];
  _RAND_28 = {2{`RANDOM}};
  mem_28 = _RAND_28[61:0];
  _RAND_29 = {2{`RANDOM}};
  mem_29 = _RAND_29[61:0];
  _RAND_30 = {2{`RANDOM}};
  mem_30 = _RAND_30[61:0];
  _RAND_31 = {2{`RANDOM}};
  mem_31 = _RAND_31[61:0];
  _RAND_32 = {2{`RANDOM}};
  mem_32 = _RAND_32[61:0];
  _RAND_33 = {2{`RANDOM}};
  mem_33 = _RAND_33[61:0];
  _RAND_34 = {2{`RANDOM}};
  mem_34 = _RAND_34[61:0];
  _RAND_35 = {2{`RANDOM}};
  mem_35 = _RAND_35[61:0];
  _RAND_36 = {2{`RANDOM}};
  mem_36 = _RAND_36[61:0];
  _RAND_37 = {2{`RANDOM}};
  mem_37 = _RAND_37[61:0];
  _RAND_38 = {2{`RANDOM}};
  mem_38 = _RAND_38[61:0];
  _RAND_39 = {2{`RANDOM}};
  mem_39 = _RAND_39[61:0];
  _RAND_40 = {2{`RANDOM}};
  mem_40 = _RAND_40[61:0];
  _RAND_41 = {2{`RANDOM}};
  mem_41 = _RAND_41[61:0];
  _RAND_42 = {2{`RANDOM}};
  mem_42 = _RAND_42[61:0];
  _RAND_43 = {2{`RANDOM}};
  mem_43 = _RAND_43[61:0];
  _RAND_44 = {2{`RANDOM}};
  mem_44 = _RAND_44[61:0];
  _RAND_45 = {2{`RANDOM}};
  mem_45 = _RAND_45[61:0];
  _RAND_46 = {2{`RANDOM}};
  mem_46 = _RAND_46[61:0];
  _RAND_47 = {2{`RANDOM}};
  mem_47 = _RAND_47[61:0];
  _RAND_48 = {2{`RANDOM}};
  mem_48 = _RAND_48[61:0];
  _RAND_49 = {2{`RANDOM}};
  mem_49 = _RAND_49[61:0];
  _RAND_50 = {2{`RANDOM}};
  mem_50 = _RAND_50[61:0];
  _RAND_51 = {2{`RANDOM}};
  mem_51 = _RAND_51[61:0];
  _RAND_52 = {2{`RANDOM}};
  mem_52 = _RAND_52[61:0];
  _RAND_53 = {2{`RANDOM}};
  mem_53 = _RAND_53[61:0];
  _RAND_54 = {2{`RANDOM}};
  mem_54 = _RAND_54[61:0];
  _RAND_55 = {2{`RANDOM}};
  mem_55 = _RAND_55[61:0];
  _RAND_56 = {2{`RANDOM}};
  mem_56 = _RAND_56[61:0];
  _RAND_57 = {2{`RANDOM}};
  mem_57 = _RAND_57[61:0];
  _RAND_58 = {2{`RANDOM}};
  mem_58 = _RAND_58[61:0];
  _RAND_59 = {2{`RANDOM}};
  mem_59 = _RAND_59[61:0];
  _RAND_60 = {2{`RANDOM}};
  mem_60 = _RAND_60[61:0];
  _RAND_61 = {2{`RANDOM}};
  mem_61 = _RAND_61[61:0];
  _RAND_62 = {2{`RANDOM}};
  mem_62 = _RAND_62[61:0];
  _RAND_63 = {2{`RANDOM}};
  mem_63 = _RAND_63[61:0];
  _RAND_64 = {2{`RANDOM}};
  mem_64 = _RAND_64[61:0];
  _RAND_65 = {2{`RANDOM}};
  mem_65 = _RAND_65[61:0];
  _RAND_66 = {2{`RANDOM}};
  mem_66 = _RAND_66[61:0];
  _RAND_67 = {2{`RANDOM}};
  mem_67 = _RAND_67[61:0];
  _RAND_68 = {2{`RANDOM}};
  mem_68 = _RAND_68[61:0];
  _RAND_69 = {2{`RANDOM}};
  mem_69 = _RAND_69[61:0];
  _RAND_70 = {2{`RANDOM}};
  mem_70 = _RAND_70[61:0];
  _RAND_71 = {2{`RANDOM}};
  mem_71 = _RAND_71[61:0];
  _RAND_72 = {2{`RANDOM}};
  mem_72 = _RAND_72[61:0];
  _RAND_73 = {2{`RANDOM}};
  mem_73 = _RAND_73[61:0];
  _RAND_74 = {2{`RANDOM}};
  mem_74 = _RAND_74[61:0];
  _RAND_75 = {2{`RANDOM}};
  mem_75 = _RAND_75[61:0];
  _RAND_76 = {2{`RANDOM}};
  mem_76 = _RAND_76[61:0];
  _RAND_77 = {2{`RANDOM}};
  mem_77 = _RAND_77[61:0];
  _RAND_78 = {2{`RANDOM}};
  mem_78 = _RAND_78[61:0];
  _RAND_79 = {2{`RANDOM}};
  mem_79 = _RAND_79[61:0];
  _RAND_80 = {2{`RANDOM}};
  mem_80 = _RAND_80[61:0];
  _RAND_81 = {2{`RANDOM}};
  mem_81 = _RAND_81[61:0];
  _RAND_82 = {2{`RANDOM}};
  mem_82 = _RAND_82[61:0];
  _RAND_83 = {2{`RANDOM}};
  mem_83 = _RAND_83[61:0];
  _RAND_84 = {2{`RANDOM}};
  mem_84 = _RAND_84[61:0];
  _RAND_85 = {2{`RANDOM}};
  mem_85 = _RAND_85[61:0];
  _RAND_86 = {2{`RANDOM}};
  mem_86 = _RAND_86[61:0];
  _RAND_87 = {2{`RANDOM}};
  mem_87 = _RAND_87[61:0];
  _RAND_88 = {2{`RANDOM}};
  mem_88 = _RAND_88[61:0];
  _RAND_89 = {2{`RANDOM}};
  mem_89 = _RAND_89[61:0];
  _RAND_90 = {2{`RANDOM}};
  mem_90 = _RAND_90[61:0];
  _RAND_91 = {2{`RANDOM}};
  mem_91 = _RAND_91[61:0];
  _RAND_92 = {2{`RANDOM}};
  mem_92 = _RAND_92[61:0];
  _RAND_93 = {2{`RANDOM}};
  mem_93 = _RAND_93[61:0];
  _RAND_94 = {2{`RANDOM}};
  mem_94 = _RAND_94[61:0];
  _RAND_95 = {2{`RANDOM}};
  mem_95 = _RAND_95[61:0];
  _RAND_96 = {2{`RANDOM}};
  mem_96 = _RAND_96[61:0];
  _RAND_97 = {2{`RANDOM}};
  mem_97 = _RAND_97[61:0];
  _RAND_98 = {2{`RANDOM}};
  mem_98 = _RAND_98[61:0];
  _RAND_99 = {2{`RANDOM}};
  mem_99 = _RAND_99[61:0];
  _RAND_100 = {2{`RANDOM}};
  mem_100 = _RAND_100[61:0];
  _RAND_101 = {2{`RANDOM}};
  mem_101 = _RAND_101[61:0];
  _RAND_102 = {2{`RANDOM}};
  mem_102 = _RAND_102[61:0];
  _RAND_103 = {2{`RANDOM}};
  mem_103 = _RAND_103[61:0];
  _RAND_104 = {2{`RANDOM}};
  mem_104 = _RAND_104[61:0];
  _RAND_105 = {2{`RANDOM}};
  mem_105 = _RAND_105[61:0];
  _RAND_106 = {2{`RANDOM}};
  mem_106 = _RAND_106[61:0];
  _RAND_107 = {2{`RANDOM}};
  mem_107 = _RAND_107[61:0];
  _RAND_108 = {2{`RANDOM}};
  mem_108 = _RAND_108[61:0];
  _RAND_109 = {2{`RANDOM}};
  mem_109 = _RAND_109[61:0];
  _RAND_110 = {2{`RANDOM}};
  mem_110 = _RAND_110[61:0];
  _RAND_111 = {2{`RANDOM}};
  mem_111 = _RAND_111[61:0];
  _RAND_112 = {2{`RANDOM}};
  mem_112 = _RAND_112[61:0];
  _RAND_113 = {2{`RANDOM}};
  mem_113 = _RAND_113[61:0];
  _RAND_114 = {2{`RANDOM}};
  mem_114 = _RAND_114[61:0];
  _RAND_115 = {2{`RANDOM}};
  mem_115 = _RAND_115[61:0];
  _RAND_116 = {2{`RANDOM}};
  mem_116 = _RAND_116[61:0];
  _RAND_117 = {2{`RANDOM}};
  mem_117 = _RAND_117[61:0];
  _RAND_118 = {2{`RANDOM}};
  mem_118 = _RAND_118[61:0];
  _RAND_119 = {2{`RANDOM}};
  mem_119 = _RAND_119[61:0];
  _RAND_120 = {2{`RANDOM}};
  mem_120 = _RAND_120[61:0];
  _RAND_121 = {2{`RANDOM}};
  mem_121 = _RAND_121[61:0];
  _RAND_122 = {2{`RANDOM}};
  mem_122 = _RAND_122[61:0];
  _RAND_123 = {2{`RANDOM}};
  mem_123 = _RAND_123[61:0];
  _RAND_124 = {2{`RANDOM}};
  mem_124 = _RAND_124[61:0];
  _RAND_125 = {2{`RANDOM}};
  mem_125 = _RAND_125[61:0];
  _RAND_126 = {2{`RANDOM}};
  mem_126 = _RAND_126[61:0];
  _RAND_127 = {2{`RANDOM}};
  mem_127 = _RAND_127[61:0];
  _RAND_128 = {2{`RANDOM}};
  mem_128 = _RAND_128[61:0];
  _RAND_129 = {2{`RANDOM}};
  mem_129 = _RAND_129[61:0];
  _RAND_130 = {2{`RANDOM}};
  mem_130 = _RAND_130[61:0];
  _RAND_131 = {2{`RANDOM}};
  mem_131 = _RAND_131[61:0];
  _RAND_132 = {2{`RANDOM}};
  mem_132 = _RAND_132[61:0];
  _RAND_133 = {2{`RANDOM}};
  mem_133 = _RAND_133[61:0];
  _RAND_134 = {2{`RANDOM}};
  mem_134 = _RAND_134[61:0];
  _RAND_135 = {2{`RANDOM}};
  mem_135 = _RAND_135[61:0];
  _RAND_136 = {2{`RANDOM}};
  mem_136 = _RAND_136[61:0];
  _RAND_137 = {2{`RANDOM}};
  mem_137 = _RAND_137[61:0];
  _RAND_138 = {2{`RANDOM}};
  mem_138 = _RAND_138[61:0];
  _RAND_139 = {2{`RANDOM}};
  mem_139 = _RAND_139[61:0];
  _RAND_140 = {2{`RANDOM}};
  mem_140 = _RAND_140[61:0];
  _RAND_141 = {2{`RANDOM}};
  mem_141 = _RAND_141[61:0];
  _RAND_142 = {2{`RANDOM}};
  mem_142 = _RAND_142[61:0];
  _RAND_143 = {2{`RANDOM}};
  mem_143 = _RAND_143[61:0];
  _RAND_144 = {2{`RANDOM}};
  mem_144 = _RAND_144[61:0];
  _RAND_145 = {2{`RANDOM}};
  mem_145 = _RAND_145[61:0];
  _RAND_146 = {2{`RANDOM}};
  mem_146 = _RAND_146[61:0];
  _RAND_147 = {2{`RANDOM}};
  mem_147 = _RAND_147[61:0];
  _RAND_148 = {2{`RANDOM}};
  mem_148 = _RAND_148[61:0];
  _RAND_149 = {2{`RANDOM}};
  mem_149 = _RAND_149[61:0];
  _RAND_150 = {2{`RANDOM}};
  mem_150 = _RAND_150[61:0];
  _RAND_151 = {2{`RANDOM}};
  mem_151 = _RAND_151[61:0];
  _RAND_152 = {2{`RANDOM}};
  mem_152 = _RAND_152[61:0];
  _RAND_153 = {2{`RANDOM}};
  mem_153 = _RAND_153[61:0];
  _RAND_154 = {2{`RANDOM}};
  mem_154 = _RAND_154[61:0];
  _RAND_155 = {2{`RANDOM}};
  mem_155 = _RAND_155[61:0];
  _RAND_156 = {2{`RANDOM}};
  mem_156 = _RAND_156[61:0];
  _RAND_157 = {2{`RANDOM}};
  mem_157 = _RAND_157[61:0];
  _RAND_158 = {2{`RANDOM}};
  mem_158 = _RAND_158[61:0];
  _RAND_159 = {2{`RANDOM}};
  mem_159 = _RAND_159[61:0];
  _RAND_160 = {2{`RANDOM}};
  mem_160 = _RAND_160[61:0];
  _RAND_161 = {2{`RANDOM}};
  mem_161 = _RAND_161[61:0];
  _RAND_162 = {2{`RANDOM}};
  mem_162 = _RAND_162[61:0];
  _RAND_163 = {2{`RANDOM}};
  mem_163 = _RAND_163[61:0];
  _RAND_164 = {2{`RANDOM}};
  mem_164 = _RAND_164[61:0];
  _RAND_165 = {2{`RANDOM}};
  mem_165 = _RAND_165[61:0];
  _RAND_166 = {2{`RANDOM}};
  mem_166 = _RAND_166[61:0];
  _RAND_167 = {2{`RANDOM}};
  mem_167 = _RAND_167[61:0];
  _RAND_168 = {2{`RANDOM}};
  mem_168 = _RAND_168[61:0];
  _RAND_169 = {2{`RANDOM}};
  mem_169 = _RAND_169[61:0];
  _RAND_170 = {2{`RANDOM}};
  mem_170 = _RAND_170[61:0];
  _RAND_171 = {2{`RANDOM}};
  mem_171 = _RAND_171[61:0];
  _RAND_172 = {2{`RANDOM}};
  mem_172 = _RAND_172[61:0];
  _RAND_173 = {2{`RANDOM}};
  mem_173 = _RAND_173[61:0];
  _RAND_174 = {2{`RANDOM}};
  mem_174 = _RAND_174[61:0];
  _RAND_175 = {2{`RANDOM}};
  mem_175 = _RAND_175[61:0];
  _RAND_176 = {2{`RANDOM}};
  mem_176 = _RAND_176[61:0];
  _RAND_177 = {2{`RANDOM}};
  mem_177 = _RAND_177[61:0];
  _RAND_178 = {2{`RANDOM}};
  mem_178 = _RAND_178[61:0];
  _RAND_179 = {2{`RANDOM}};
  mem_179 = _RAND_179[61:0];
  _RAND_180 = {2{`RANDOM}};
  mem_180 = _RAND_180[61:0];
  _RAND_181 = {2{`RANDOM}};
  mem_181 = _RAND_181[61:0];
  _RAND_182 = {2{`RANDOM}};
  mem_182 = _RAND_182[61:0];
  _RAND_183 = {2{`RANDOM}};
  mem_183 = _RAND_183[61:0];
  _RAND_184 = {2{`RANDOM}};
  mem_184 = _RAND_184[61:0];
  _RAND_185 = {2{`RANDOM}};
  mem_185 = _RAND_185[61:0];
  _RAND_186 = {2{`RANDOM}};
  mem_186 = _RAND_186[61:0];
  _RAND_187 = {2{`RANDOM}};
  mem_187 = _RAND_187[61:0];
  _RAND_188 = {2{`RANDOM}};
  mem_188 = _RAND_188[61:0];
  _RAND_189 = {2{`RANDOM}};
  mem_189 = _RAND_189[61:0];
  _RAND_190 = {2{`RANDOM}};
  mem_190 = _RAND_190[61:0];
  _RAND_191 = {2{`RANDOM}};
  mem_191 = _RAND_191[61:0];
  _RAND_192 = {2{`RANDOM}};
  mem_192 = _RAND_192[61:0];
  _RAND_193 = {2{`RANDOM}};
  mem_193 = _RAND_193[61:0];
  _RAND_194 = {2{`RANDOM}};
  mem_194 = _RAND_194[61:0];
  _RAND_195 = {2{`RANDOM}};
  mem_195 = _RAND_195[61:0];
  _RAND_196 = {2{`RANDOM}};
  mem_196 = _RAND_196[61:0];
  _RAND_197 = {2{`RANDOM}};
  mem_197 = _RAND_197[61:0];
  _RAND_198 = {2{`RANDOM}};
  mem_198 = _RAND_198[61:0];
  _RAND_199 = {2{`RANDOM}};
  mem_199 = _RAND_199[61:0];
  _RAND_200 = {2{`RANDOM}};
  mem_200 = _RAND_200[61:0];
  _RAND_201 = {2{`RANDOM}};
  mem_201 = _RAND_201[61:0];
  _RAND_202 = {2{`RANDOM}};
  mem_202 = _RAND_202[61:0];
  _RAND_203 = {2{`RANDOM}};
  mem_203 = _RAND_203[61:0];
  _RAND_204 = {2{`RANDOM}};
  mem_204 = _RAND_204[61:0];
  _RAND_205 = {2{`RANDOM}};
  mem_205 = _RAND_205[61:0];
  _RAND_206 = {2{`RANDOM}};
  mem_206 = _RAND_206[61:0];
  _RAND_207 = {2{`RANDOM}};
  mem_207 = _RAND_207[61:0];
  _RAND_208 = {2{`RANDOM}};
  mem_208 = _RAND_208[61:0];
  _RAND_209 = {2{`RANDOM}};
  mem_209 = _RAND_209[61:0];
  _RAND_210 = {2{`RANDOM}};
  mem_210 = _RAND_210[61:0];
  _RAND_211 = {2{`RANDOM}};
  mem_211 = _RAND_211[61:0];
  _RAND_212 = {2{`RANDOM}};
  mem_212 = _RAND_212[61:0];
  _RAND_213 = {2{`RANDOM}};
  mem_213 = _RAND_213[61:0];
  _RAND_214 = {2{`RANDOM}};
  mem_214 = _RAND_214[61:0];
  _RAND_215 = {2{`RANDOM}};
  mem_215 = _RAND_215[61:0];
  _RAND_216 = {2{`RANDOM}};
  mem_216 = _RAND_216[61:0];
  _RAND_217 = {2{`RANDOM}};
  mem_217 = _RAND_217[61:0];
  _RAND_218 = {2{`RANDOM}};
  mem_218 = _RAND_218[61:0];
  _RAND_219 = {2{`RANDOM}};
  mem_219 = _RAND_219[61:0];
  _RAND_220 = {2{`RANDOM}};
  mem_220 = _RAND_220[61:0];
  _RAND_221 = {2{`RANDOM}};
  mem_221 = _RAND_221[61:0];
  _RAND_222 = {2{`RANDOM}};
  mem_222 = _RAND_222[61:0];
  _RAND_223 = {2{`RANDOM}};
  mem_223 = _RAND_223[61:0];
  _RAND_224 = {2{`RANDOM}};
  mem_224 = _RAND_224[61:0];
  _RAND_225 = {2{`RANDOM}};
  mem_225 = _RAND_225[61:0];
  _RAND_226 = {2{`RANDOM}};
  mem_226 = _RAND_226[61:0];
  _RAND_227 = {2{`RANDOM}};
  mem_227 = _RAND_227[61:0];
  _RAND_228 = {2{`RANDOM}};
  mem_228 = _RAND_228[61:0];
  _RAND_229 = {2{`RANDOM}};
  mem_229 = _RAND_229[61:0];
  _RAND_230 = {2{`RANDOM}};
  mem_230 = _RAND_230[61:0];
  _RAND_231 = {2{`RANDOM}};
  mem_231 = _RAND_231[61:0];
  _RAND_232 = {2{`RANDOM}};
  mem_232 = _RAND_232[61:0];
  _RAND_233 = {2{`RANDOM}};
  mem_233 = _RAND_233[61:0];
  _RAND_234 = {2{`RANDOM}};
  mem_234 = _RAND_234[61:0];
  _RAND_235 = {2{`RANDOM}};
  mem_235 = _RAND_235[61:0];
  _RAND_236 = {2{`RANDOM}};
  mem_236 = _RAND_236[61:0];
  _RAND_237 = {2{`RANDOM}};
  mem_237 = _RAND_237[61:0];
  _RAND_238 = {2{`RANDOM}};
  mem_238 = _RAND_238[61:0];
  _RAND_239 = {2{`RANDOM}};
  mem_239 = _RAND_239[61:0];
  _RAND_240 = {2{`RANDOM}};
  mem_240 = _RAND_240[61:0];
  _RAND_241 = {2{`RANDOM}};
  mem_241 = _RAND_241[61:0];
  _RAND_242 = {2{`RANDOM}};
  mem_242 = _RAND_242[61:0];
  _RAND_243 = {2{`RANDOM}};
  mem_243 = _RAND_243[61:0];
  _RAND_244 = {2{`RANDOM}};
  mem_244 = _RAND_244[61:0];
  _RAND_245 = {2{`RANDOM}};
  mem_245 = _RAND_245[61:0];
  _RAND_246 = {2{`RANDOM}};
  mem_246 = _RAND_246[61:0];
  _RAND_247 = {2{`RANDOM}};
  mem_247 = _RAND_247[61:0];
  _RAND_248 = {2{`RANDOM}};
  mem_248 = _RAND_248[61:0];
  _RAND_249 = {2{`RANDOM}};
  mem_249 = _RAND_249[61:0];
  _RAND_250 = {2{`RANDOM}};
  mem_250 = _RAND_250[61:0];
  _RAND_251 = {2{`RANDOM}};
  mem_251 = _RAND_251[61:0];
  _RAND_252 = {2{`RANDOM}};
  mem_252 = _RAND_252[61:0];
  _RAND_253 = {2{`RANDOM}};
  mem_253 = _RAND_253[61:0];
  _RAND_254 = {2{`RANDOM}};
  mem_254 = _RAND_254[61:0];
  _RAND_255 = {2{`RANDOM}};
  mem_255 = _RAND_255[61:0];
  _RAND_256 = {2{`RANDOM}};
  io_douta_REG = _RAND_256[61:0];
  _RAND_257 = {2{`RANDOM}};
  io_doutb_REG = _RAND_257[61:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM_1(
  input         clock,
  input         reset,
  input         io_wea,
  input  [7:0]  io_addra,
  input  [7:0]  io_addrb,
  input  [61:0] io_dina,
  output [61:0] io_douta,
  output [61:0] io_doutb
);
  wire  sim_dual_port_bram_clock; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_reset; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_io_wea; // @[RAMWrapper.scala 30:36]
  wire [7:0] sim_dual_port_bram_io_addra; // @[RAMWrapper.scala 30:36]
  wire [7:0] sim_dual_port_bram_io_addrb; // @[RAMWrapper.scala 30:36]
  wire [61:0] sim_dual_port_bram_io_dina; // @[RAMWrapper.scala 30:36]
  wire [61:0] sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 30:36]
  wire [61:0] sim_dual_port_bram_io_doutb; // @[RAMWrapper.scala 30:36]
  SimDualPortBRAM_1 sim_dual_port_bram ( // @[RAMWrapper.scala 30:36]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_wea(sim_dual_port_bram_io_wea),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dina(sim_dual_port_bram_io_dina),
    .io_douta(sim_dual_port_bram_io_douta),
    .io_doutb(sim_dual_port_bram_io_doutb)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 31:27]
  assign io_doutb = sim_dual_port_bram_io_doutb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_wea = io_wea; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_dina = io_dina; // @[RAMWrapper.scala 31:27]
endmodule
module BPU(
  input         clock,
  input         reset,
  input  [63:0] io_req_next_line,
  output        io_resp_taken_vec_0,
  output        io_resp_taken_vec_1,
  output [63:0] io_resp_target_0,
  output [63:0] io_resp_target_1,
  input         io_update_dec_v,
  input  [63:0] io_update_dec_pc_br,
  input         io_update_exe_v,
  input         io_update_exe_errpr,
  input  [63:0] io_update_exe_pc_br,
  input  [63:0] io_update_exe_target,
  input         io_update_exe_taken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  history_clock; // @[BPU.scala 86:23]
  wire  history_reset; // @[BPU.scala 86:23]
  wire  history_io_wea; // @[BPU.scala 86:23]
  wire [7:0] history_io_addra; // @[BPU.scala 86:23]
  wire [7:0] history_io_addrb; // @[BPU.scala 86:23]
  wire [1:0] history_io_dina; // @[BPU.scala 86:23]
  wire [1:0] history_io_douta; // @[BPU.scala 86:23]
  wire [1:0] history_io_doutb; // @[BPU.scala 86:23]
  wire  buffer_clock; // @[BPU.scala 87:23]
  wire  buffer_reset; // @[BPU.scala 87:23]
  wire  buffer_io_wea; // @[BPU.scala 87:23]
  wire [7:0] buffer_io_addra; // @[BPU.scala 87:23]
  wire [7:0] buffer_io_addrb; // @[BPU.scala 87:23]
  wire [61:0] buffer_io_dina; // @[BPU.scala 87:23]
  wire [61:0] buffer_io_douta; // @[BPU.scala 87:23]
  wire [61:0] buffer_io_doutb; // @[BPU.scala 87:23]
  reg [7:0] bht_cache_tag_0; // @[BPU.scala 77:27]
  reg [1:0] bht_cache_stat_0; // @[BPU.scala 78:31]
  reg  cache_or_update_hit; // @[BPU.scala 82:32]
  reg [1:0] chosen_result; // @[BPU.scala 83:26]
  wire  _waddr_T = ~io_update_dec_v; // @[BPU.scala 90:24]
  wire [63:0] waddr = ~io_update_dec_v ? io_update_exe_pc_br : io_update_dec_pc_br; // @[BPU.scala 90:23]
  wire  exe_update = io_update_exe_taken ? ~(&io_update_exe_pc_br[1:0]) : |io_update_exe_pc_br[1:0]; // @[BPU.scala 91:23]
  wire  _update_T_2 = ~io_update_exe_v ? 1'h0 : exe_update; // @[BPU.scala 92:45]
  wire  update = _waddr_T ? _update_T_2 : 1'h1; // @[BPU.scala 92:23]
  wire [1:0] _wdata_T_3 = io_update_exe_pc_br[1:0] + 2'h1; // @[BPU.scala 93:93]
  wire [1:0] _wdata_T_6 = io_update_exe_pc_br[1:0] - 2'h1; // @[BPU.scala 93:126]
  wire [1:0] _wdata_T_7 = io_update_exe_taken ? _wdata_T_3 : _wdata_T_6; // @[BPU.scala 93:45]
  wire [1:0] _wdata_T_10 = io_update_dec_pc_br[1:0] - 2'h1; // @[BPU.scala 93:160]
  wire  history_io_addra_higher_hi_hi_hi = waddr[16] ^ waddr[15] ^ waddr[9]; // @[BPU.scala 60:56]
  wire  history_io_addra_higher_hi_hi_lo = waddr[15] ^ waddr[14] ^ waddr[8]; // @[BPU.scala 60:105]
  wire  history_io_addra_higher_hi_lo = waddr[14] ^ waddr[13] ^ waddr[7]; // @[BPU.scala 60:154]
  wire  history_io_addra_higher_lo_hi_hi = waddr[13] ^ waddr[12] ^ waddr[6]; // @[BPU.scala 60:203]
  wire  history_io_addra_higher_lo_hi_lo = waddr[12] ^ waddr[11] ^ waddr[5]; // @[BPU.scala 60:252]
  wire  history_io_addra_higher_lo_lo = waddr[11] ^ waddr[10] ^ waddr[4]; // @[BPU.scala 60:300]
  wire  history_io_addra_lo = waddr[10] ^ waddr[9] ^ waddr[3]; // @[BPU.scala 64:40]
  wire  history_io_addra_lo_1 = waddr[2]; // @[BPU.scala 74:35]
  wire [7:0] _history_io_addra_T_4 = {history_io_addra_higher_hi_hi_hi,history_io_addra_higher_hi_hi_lo,
    history_io_addra_higher_hi_lo,history_io_addra_higher_lo_hi_hi,history_io_addra_higher_lo_hi_lo,
    history_io_addra_higher_lo_lo,history_io_addra_lo,history_io_addra_lo_1}; // @[Cat.scala 30:58]
  wire  history_io_addra_higher_hi_hi_hi_1 = io_req_next_line[16] ^ io_req_next_line[15] ^ io_req_next_line[9]; // @[BPU.scala 60:56]
  wire  history_io_addra_higher_hi_hi_lo_1 = io_req_next_line[15] ^ io_req_next_line[14] ^ io_req_next_line[8]; // @[BPU.scala 60:105]
  wire  history_io_addra_higher_hi_lo_1 = io_req_next_line[14] ^ io_req_next_line[13] ^ io_req_next_line[7]; // @[BPU.scala 60:154]
  wire  history_io_addra_higher_lo_hi_hi_1 = io_req_next_line[13] ^ io_req_next_line[12] ^ io_req_next_line[6]; // @[BPU.scala 60:203]
  wire  history_io_addra_higher_lo_hi_lo_1 = io_req_next_line[12] ^ io_req_next_line[11] ^ io_req_next_line[5]; // @[BPU.scala 60:252]
  wire  history_io_addra_higher_lo_lo_1 = io_req_next_line[11] ^ io_req_next_line[10] ^ io_req_next_line[4]; // @[BPU.scala 60:300]
  wire  history_io_addra_lo_2 = io_req_next_line[10] ^ io_req_next_line[9] ^ io_req_next_line[3]; // @[BPU.scala 64:40]
  wire [6:0] history_io_addra_hi_3 = {history_io_addra_higher_hi_hi_hi_1,history_io_addra_higher_hi_hi_lo_1,
    history_io_addra_higher_hi_lo_1,history_io_addra_higher_lo_hi_hi_1,history_io_addra_higher_lo_hi_lo_1,
    history_io_addra_higher_lo_lo_1,history_io_addra_lo_2}; // @[Cat.scala 30:58]
  wire  history_io_addra_lo_3 = io_req_next_line[2]; // @[BPU.scala 74:35]
  wire [7:0] _history_io_addra_T_9 = {history_io_addra_higher_hi_hi_hi_1,history_io_addra_higher_hi_hi_lo_1,
    history_io_addra_higher_hi_lo_1,history_io_addra_higher_lo_hi_hi_1,history_io_addra_higher_lo_hi_lo_1,
    history_io_addra_higher_lo_lo_1,history_io_addra_lo_2,history_io_addra_lo_3}; // @[Cat.scala 30:58]
  wire [63:0] _history_io_addrb_T_1 = io_req_next_line + 64'h4; // @[BPU.scala 98:60]
  wire  history_io_addrb_higher_hi_hi_hi = _history_io_addrb_T_1[16] ^ _history_io_addrb_T_1[15] ^ _history_io_addrb_T_1
    [9]; // @[BPU.scala 60:56]
  wire  history_io_addrb_higher_hi_hi_lo = _history_io_addrb_T_1[15] ^ _history_io_addrb_T_1[14] ^ _history_io_addrb_T_1
    [8]; // @[BPU.scala 60:105]
  wire  history_io_addrb_higher_hi_lo = _history_io_addrb_T_1[14] ^ _history_io_addrb_T_1[13] ^ _history_io_addrb_T_1[7]
    ; // @[BPU.scala 60:154]
  wire  history_io_addrb_higher_lo_hi_hi = _history_io_addrb_T_1[13] ^ _history_io_addrb_T_1[12] ^ _history_io_addrb_T_1
    [6]; // @[BPU.scala 60:203]
  wire  history_io_addrb_higher_lo_hi_lo = _history_io_addrb_T_1[12] ^ _history_io_addrb_T_1[11] ^ _history_io_addrb_T_1
    [5]; // @[BPU.scala 60:252]
  wire  history_io_addrb_higher_lo_lo = _history_io_addrb_T_1[11] ^ _history_io_addrb_T_1[10] ^ _history_io_addrb_T_1[4]
    ; // @[BPU.scala 60:300]
  wire  history_io_addrb_lo = _history_io_addrb_T_1[10] ^ _history_io_addrb_T_1[9] ^ _history_io_addrb_T_1[3]; // @[BPU.scala 64:40]
  wire [6:0] history_io_addrb_hi_1 = {history_io_addrb_higher_hi_hi_hi,history_io_addrb_higher_hi_hi_lo,
    history_io_addrb_higher_hi_lo,history_io_addrb_higher_lo_hi_hi,history_io_addrb_higher_lo_hi_lo,
    history_io_addrb_higher_lo_lo,history_io_addrb_lo}; // @[Cat.scala 30:58]
  wire  history_io_addrb_lo_1 = _history_io_addrb_T_1[2]; // @[BPU.scala 74:35]
  reg  last_update; // @[BPU.scala 104:28]
  wire [1:0] _bht_first_T_1 = cache_or_update_hit ? chosen_result : 2'h0; // @[BPU.scala 105:41]
  wire [1:0] bht_first = last_update ? _bht_first_T_1 : history_io_douta; // @[BPU.scala 105:24]
  wire [63:0] _buffer_io_addra_T = io_update_exe_errpr ? io_update_exe_pc_br : io_req_next_line; // @[BPU.scala 115:45]
  wire  buffer_io_addra_higher_hi_hi_hi = _buffer_io_addra_T[16] ^ _buffer_io_addra_T[15] ^ _buffer_io_addra_T[9]; // @[BPU.scala 60:56]
  wire  buffer_io_addra_higher_hi_hi_lo = _buffer_io_addra_T[15] ^ _buffer_io_addra_T[14] ^ _buffer_io_addra_T[8]; // @[BPU.scala 60:105]
  wire  buffer_io_addra_higher_hi_lo = _buffer_io_addra_T[14] ^ _buffer_io_addra_T[13] ^ _buffer_io_addra_T[7]; // @[BPU.scala 60:154]
  wire  buffer_io_addra_higher_lo_hi_hi = _buffer_io_addra_T[13] ^ _buffer_io_addra_T[12] ^ _buffer_io_addra_T[6]; // @[BPU.scala 60:203]
  wire  buffer_io_addra_higher_lo_hi_lo = _buffer_io_addra_T[12] ^ _buffer_io_addra_T[11] ^ _buffer_io_addra_T[5]; // @[BPU.scala 60:252]
  wire  buffer_io_addra_higher_lo_lo = _buffer_io_addra_T[11] ^ _buffer_io_addra_T[10] ^ _buffer_io_addra_T[4]; // @[BPU.scala 60:300]
  wire  buffer_io_addra_lo = _buffer_io_addra_T[10] ^ _buffer_io_addra_T[9] ^ _buffer_io_addra_T[3]; // @[BPU.scala 64:40]
  wire [6:0] buffer_io_addra_hi_1 = {buffer_io_addra_higher_hi_hi_hi,buffer_io_addra_higher_hi_hi_lo,
    buffer_io_addra_higher_hi_lo,buffer_io_addra_higher_lo_hi_hi,buffer_io_addra_higher_lo_hi_lo,
    buffer_io_addra_higher_lo_lo,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  wire  buffer_io_addra_lo_1 = _buffer_io_addra_T[2]; // @[BPU.scala 74:35]
  reg  io_resp_target_0_REG; // @[BPU.scala 121:39]
  reg [61:0] io_resp_target_0_REG_1; // @[BPU.scala 121:63]
  wire [61:0] io_resp_target_0_hi = io_resp_target_0_REG ? io_resp_target_0_REG_1 : buffer_io_douta; // @[BPU.scala 121:31]
  wire  hit_in_bht_cache = bht_cache_tag_0 == _history_io_addra_T_9; // @[BPU.scala 128:28]
  reg [7:0] bht_cache_tag_0_REG; // @[BPU.scala 143:49]
  wire  update_query_hit = _history_io_addra_T_9 == _history_io_addra_T_4; // @[BPU.scala 148:64]
  DualPortBRAM history ( // @[BPU.scala 86:23]
    .clock(history_clock),
    .reset(history_reset),
    .io_wea(history_io_wea),
    .io_addra(history_io_addra),
    .io_addrb(history_io_addrb),
    .io_dina(history_io_dina),
    .io_douta(history_io_douta),
    .io_doutb(history_io_doutb)
  );
  DualPortBRAM_1 buffer ( // @[BPU.scala 87:23]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .io_wea(buffer_io_wea),
    .io_addra(buffer_io_addra),
    .io_addrb(buffer_io_addrb),
    .io_dina(buffer_io_dina),
    .io_douta(buffer_io_douta),
    .io_doutb(buffer_io_doutb)
  );
  assign io_resp_taken_vec_0 = bht_first[1]; // @[BPU.scala 107:36]
  assign io_resp_taken_vec_1 = history_io_doutb[1]; // @[BPU.scala 108:43]
  assign io_resp_target_0 = {io_resp_target_0_hi,bht_first}; // @[Cat.scala 30:58]
  assign io_resp_target_1 = {buffer_io_doutb,history_io_doutb}; // @[Cat.scala 30:58]
  assign history_clock = clock;
  assign history_reset = reset;
  assign history_io_wea = _waddr_T ? _update_T_2 : 1'h1; // @[BPU.scala 92:23]
  assign history_io_addra = update ? _history_io_addra_T_4 : _history_io_addra_T_9; // @[BPU.scala 97:26]
  assign history_io_addrb = {history_io_addrb_hi_1,history_io_addrb_lo_1}; // @[Cat.scala 30:58]
  assign history_io_dina = _waddr_T ? _wdata_T_7 : _wdata_T_10; // @[BPU.scala 93:23]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_io_wea = io_update_exe_errpr & io_update_exe_v; // @[BPU.scala 113:40]
  assign buffer_io_addra = {buffer_io_addra_hi_1,buffer_io_addra_lo_1}; // @[Cat.scala 30:58]
  assign buffer_io_addrb = {history_io_addrb_hi_1,history_io_addrb_lo_1}; // @[Cat.scala 30:58]
  assign buffer_io_dina = io_update_exe_target[63:2]; // @[BPU.scala 117:41]
  always @(posedge clock) begin
    if (!(update & hit_in_bht_cache)) begin // @[BPU.scala 135:36]
      if (io_resp_taken_vec_0 & ~hit_in_bht_cache) begin // @[BPU.scala 139:57]
        bht_cache_tag_0 <= bht_cache_tag_0_REG; // @[BPU.scala 143:39]
      end
    end
    if (reset) begin // @[BPU.scala 78:31]
      bht_cache_stat_0 <= 2'h0; // @[BPU.scala 78:31]
    end else if (update & hit_in_bht_cache) begin // @[BPU.scala 135:36]
      bht_cache_stat_0 <= 2'h0; // @[BPU.scala 137:25]
    end else if (io_resp_taken_vec_0 & ~hit_in_bht_cache) begin // @[BPU.scala 139:57]
      if (last_update) begin // @[BPU.scala 105:24]
        bht_cache_stat_0 <= _bht_first_T_1;
      end else begin
        bht_cache_stat_0 <= history_io_douta;
      end
    end
    cache_or_update_hit <= hit_in_bht_cache | update_query_hit; // @[BPU.scala 149:43]
    if (update_query_hit) begin // @[BPU.scala 150:23]
      if (_waddr_T) begin // @[BPU.scala 93:23]
        if (io_update_exe_taken) begin // @[BPU.scala 93:45]
          chosen_result <= _wdata_T_3;
        end else begin
          chosen_result <= _wdata_T_6;
        end
      end else begin
        chosen_result <= _wdata_T_10;
      end
    end else begin
      chosen_result <= bht_cache_stat_0;
    end
    if (_waddr_T) begin // @[BPU.scala 92:23]
      if (~io_update_exe_v) begin // @[BPU.scala 92:45]
        last_update <= 1'h0;
      end else if (io_update_exe_taken) begin // @[BPU.scala 91:23]
        last_update <= ~(&io_update_exe_pc_br[1:0]);
      end else begin
        last_update <= |io_update_exe_pc_br[1:0];
      end
    end else begin
      last_update <= 1'h1;
    end
    io_resp_target_0_REG <= buffer_io_wea; // @[BPU.scala 121:39]
    io_resp_target_0_REG_1 <= buffer_io_dina; // @[BPU.scala 121:63]
    bht_cache_tag_0_REG <= {history_io_addra_hi_3,history_io_addra_lo_3}; // @[Cat.scala 30:58]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_cache_tag_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  bht_cache_stat_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  cache_or_update_hit = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  chosen_result = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  last_update = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_resp_target_0_REG = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  io_resp_target_0_REG_1 = _RAND_6[61:0];
  _RAND_7 = {1{`RANDOM}};
  bht_cache_tag_0_REG = _RAND_7[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PCGen(
  input         clock,
  input         reset,
  input         io_please_wait,
  input         io_redirect,
  input  [31:0] io_redirect_pc,
  output [31:0] io_pc_o,
  output        io_predict_taken_o_0,
  output        io_predict_taken_o_1,
  output [31:0] io_predict_target_o_0,
  output [31:0] io_predict_target_o_1,
  output        io_fetch_word_o,
  input         io_bpu_update_dec_v,
  input  [31:0] io_bpu_update_dec_pc_br,
  input         io_bpu_update_exe_v,
  input         io_bpu_update_exe_errpr,
  input  [31:0] io_bpu_update_exe_pc_br,
  input  [31:0] io_bpu_update_exe_target,
  input         io_bpu_update_exe_taken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  bpu_clock; // @[Frontend.scala 31:19]
  wire  bpu_reset; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_req_next_line; // @[Frontend.scala 31:19]
  wire  bpu_io_resp_taken_vec_0; // @[Frontend.scala 31:19]
  wire  bpu_io_resp_taken_vec_1; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_resp_target_0; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_resp_target_1; // @[Frontend.scala 31:19]
  wire  bpu_io_update_dec_v; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_update_dec_pc_br; // @[Frontend.scala 31:19]
  wire  bpu_io_update_exe_v; // @[Frontend.scala 31:19]
  wire  bpu_io_update_exe_errpr; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_update_exe_pc_br; // @[Frontend.scala 31:19]
  wire [63:0] bpu_io_update_exe_target; // @[Frontend.scala 31:19]
  wire  bpu_io_update_exe_taken; // @[Frontend.scala 31:19]
  reg [31:0] pc; // @[Frontend.scala 29:20]
  wire  cross_line = pc[4:2] == 3'h7; // @[Frontend.scala 33:44]
  wire [61:0] branch_target_0_hi = bpu_io_resp_target_0[63:2]; // @[Frontend.scala 36:50]
  wire [63:0] branch_target_0 = {branch_target_0_hi,2'h0}; // @[Cat.scala 30:58]
  wire [61:0] branch_target_1_hi = bpu_io_resp_target_1[63:2]; // @[Frontend.scala 36:50]
  wire [63:0] branch_target_1 = {branch_target_1_hi,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _first_target_T_1 = pc + 32'h4; // @[Frontend.scala 37:73]
  wire [63:0] first_target = bpu_io_resp_taken_vec_0 ? branch_target_0 : {{32'd0}, _first_target_T_1}; // @[Frontend.scala 37:25]
  wire [31:0] _legal_target_T_1 = pc + 32'h8; // @[Frontend.scala 41:64]
  wire [63:0] _legal_target_T_2 = bpu_io_resp_taken_vec_1 ? branch_target_1 : {{32'd0}, _legal_target_T_1}; // @[Frontend.scala 41:16]
  wire [63:0] _legal_target_T_3 = bpu_io_resp_taken_vec_0 ? branch_target_0 : _legal_target_T_2; // @[Frontend.scala 40:14]
  wire [63:0] legal_target = cross_line ? first_target : _legal_target_T_3; // @[Frontend.scala 39:13]
  wire [63:0] _npc_T = io_please_wait ? {{32'd0}, pc} : legal_target; // @[Frontend.scala 42:49]
  wire [63:0] npc = io_redirect ? {{32'd0}, io_redirect_pc} : _npc_T; // @[Frontend.scala 42:16]
  BPU bpu ( // @[Frontend.scala 31:19]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_req_next_line(bpu_io_req_next_line),
    .io_resp_taken_vec_0(bpu_io_resp_taken_vec_0),
    .io_resp_taken_vec_1(bpu_io_resp_taken_vec_1),
    .io_resp_target_0(bpu_io_resp_target_0),
    .io_resp_target_1(bpu_io_resp_target_1),
    .io_update_dec_v(bpu_io_update_dec_v),
    .io_update_dec_pc_br(bpu_io_update_dec_pc_br),
    .io_update_exe_v(bpu_io_update_exe_v),
    .io_update_exe_errpr(bpu_io_update_exe_errpr),
    .io_update_exe_pc_br(bpu_io_update_exe_pc_br),
    .io_update_exe_target(bpu_io_update_exe_target),
    .io_update_exe_taken(bpu_io_update_exe_taken)
  );
  assign io_pc_o = pc; // @[Frontend.scala 51:11]
  assign io_predict_taken_o_0 = bpu_io_resp_taken_vec_0; // @[Frontend.scala 49:23]
  assign io_predict_taken_o_1 = bpu_io_resp_taken_vec_1; // @[Frontend.scala 49:23]
  assign io_predict_target_o_0 = bpu_io_resp_target_0[31:0]; // @[Frontend.scala 50:23]
  assign io_predict_target_o_1 = bpu_io_resp_target_1[31:0]; // @[Frontend.scala 50:23]
  assign io_fetch_word_o = pc[4:2] == 3'h7; // @[Frontend.scala 33:44]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_req_next_line = io_redirect ? {{32'd0}, io_redirect_pc} : _npc_T; // @[Frontend.scala 42:16]
  assign bpu_io_update_dec_v = io_bpu_update_dec_v; // @[Frontend.scala 46:24]
  assign bpu_io_update_dec_pc_br = {{32'd0}, io_bpu_update_dec_pc_br}; // @[Frontend.scala 46:24]
  assign bpu_io_update_exe_v = io_bpu_update_exe_v; // @[Frontend.scala 46:24]
  assign bpu_io_update_exe_errpr = io_bpu_update_exe_errpr; // @[Frontend.scala 46:24]
  assign bpu_io_update_exe_pc_br = {{32'd0}, io_bpu_update_exe_pc_br}; // @[Frontend.scala 46:24]
  assign bpu_io_update_exe_target = {{32'd0}, io_bpu_update_exe_target}; // @[Frontend.scala 46:24]
  assign bpu_io_update_exe_taken = io_bpu_update_exe_taken; // @[Frontend.scala 46:24]
  always @(posedge clock) begin
    if (reset) begin // @[Frontend.scala 29:20]
      pc <= 32'h80000000; // @[Frontend.scala 29:20]
    end else begin
      pc <= npc[31:0]; // @[Frontend.scala 48:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Dec32(
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_bht_predict_taken,
  input  [31:0] io_target_pc,
  output        io_mops_illegal,
  output [3:0]  io_mops_next_pc,
  output [1:0]  io_mops_alu_mdu_lsu,
  output [3:0]  io_mops_branch_type,
  output [1:0]  io_mops_src_a,
  output [1:0]  io_mops_src_b,
  output        io_mops_write_dest,
  output [4:0]  io_mops_alu_op,
  output        io_mops_alu_expand,
  output [2:0]  io_mops_mem_width,
  output [1:0]  io_mops_write_src,
  output [4:0]  io_mops_rs1,
  output [4:0]  io_mops_rs2,
  output [4:0]  io_mops_rd,
  output [19:0] io_mops_imm,
  output [31:0] io_mops_pc,
  output        io_mops_predict_taken,
  output [31:0] io_mops_target_pc,
  output        io_mops_ysyx_debug,
  output        io_mops_ysyx_print,
  output [31:0] io_mops_inst
);
  wire [4:0] IRT = io_inst[24:20]; // @[Decode.scala 66:22]
  wire [4:0] IRS = io_inst[19:15]; // @[Decode.scala 67:22]
  wire [4:0] IRD = io_inst[11:7]; // @[Decode.scala 68:22]
  wire [11:0] CSR = io_inst[31:20]; // @[Decode.scala 69:22]
  wire [7:0] aluIIMM_hi = io_inst[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [19:0] aluIIMM = {aluIIMM_hi,CSR}; // @[Cat.scala 30:58]
  wire [19:0] aluUIMM = io_inst[31:12]; // @[Decode.scala 73:25]
  wire [5:0] shamtIMM_lo = io_inst[25:20]; // @[Decode.scala 74:52]
  wire [19:0] shamtIMM = {14'h0,shamtIMM_lo}; // @[Cat.scala 30:58]
  wire [6:0] lsuSIMM_hi_lo = io_inst[31:25]; // @[Decode.scala 76:63]
  wire [19:0] lsuSIMM = {aluIIMM_hi,lsuSIMM_hi_lo,IRD}; // @[Cat.scala 30:58]
  wire [7:0] JIMM_hi_lo = io_inst[19:12]; // @[Decode.scala 77:42]
  wire  JIMM_lo_hi = io_inst[20]; // @[Decode.scala 77:59]
  wire [9:0] JIMM_lo_lo = io_inst[30:21]; // @[Decode.scala 77:72]
  wire [19:0] JIMM = {io_inst[31],JIMM_hi_lo,JIMM_lo_hi,JIMM_lo_lo}; // @[Cat.scala 30:58]
  wire [6:0] BIMM_hi_hi_hi = io_inst[31] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire  BIMM_hi_lo = io_inst[7]; // @[Decode.scala 79:76]
  wire [5:0] BIMM_lo_hi_hi = io_inst[30:25]; // @[Decode.scala 79:88]
  wire [3:0] BIMM_lo_hi_lo = io_inst[11:8]; // @[Decode.scala 79:105]
  wire [19:0] BIMM = {BIMM_hi_hi_hi,io_inst[31],BIMM_hi_lo,BIMM_lo_hi_hi,BIMM_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] CSRIMM = {8'h0,CSR}; // @[Cat.scala 30:58]
  wire [31:0] _control_signal_T = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _control_signal_T_1 = 32'h37 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_3 = 32'h17 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_5 = 32'h6f == _control_signal_T; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_6 = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _control_signal_T_7 = 32'h67 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_9 = 32'h63 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_11 = 32'h1063 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_13 = 32'h4063 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_15 = 32'h5063 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_17 = 32'h6063 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_19 = 32'h7063 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_21 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _control_signal_T_23 = 32'h3 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_25 = 32'h1003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_27 = 32'h2003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_29 = 32'h4003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_31 = 32'h5003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_33 = 32'h23 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_35 = 32'h1023 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_37 = 32'h2023 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_39 = 32'h13 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_41 = 32'h2013 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_43 = 32'h3013 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_45 = 32'h4013 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_47 = 32'h6013 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_49 = 32'h7013 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_51 = 32'h30200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _control_signal_T_53 = 32'h10200073 == io_inst; // @[Lookup.scala 31:38]
  wire  _control_signal_T_55 = 32'h200073 == io_inst; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_56 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _control_signal_T_57 = 32'h33 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_59 = 32'h40000033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_61 = 32'h1033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_63 = 32'h2033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_65 = 32'h3033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_67 = 32'h4033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_69 = 32'h5033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_71 = 32'h40005033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_73 = 32'h6033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_75 = 32'h7033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_76 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _control_signal_T_77 = 32'h1013 == _control_signal_T_76; // @[Lookup.scala 31:38]
  wire  _control_signal_T_79 = 32'h5013 == _control_signal_T_76; // @[Lookup.scala 31:38]
  wire  _control_signal_T_81 = 32'h40005013 == _control_signal_T_76; // @[Lookup.scala 31:38]
  wire  _control_signal_T_83 = 32'h1b == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_85 = 32'h101b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_87 = 32'h501b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_89 = 32'h4000501b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_91 = 32'h3b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_93 = 32'h4000003b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_95 = 32'h103b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_97 = 32'h503b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_99 = 32'h4000503b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_101 = 32'h3003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_103 = 32'h6003 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_105 = 32'h3023 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_107 = 32'h2000033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_109 = 32'h2001033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_111 = 32'h2002033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_113 = 32'h2003033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_115 = 32'h2004033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_117 = 32'h2005033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_119 = 32'h2006033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_121 = 32'h2007033 == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_123 = 32'h200003b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_125 = 32'h200403b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_127 = 32'h200503b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_129 = 32'h200603b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_131 = 32'h200703b == _control_signal_T_56; // @[Lookup.scala 31:38]
  wire  _control_signal_T_133 = 32'h1073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_135 = 32'h2073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_137 = 32'h3073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_139 = 32'h5073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_141 = 32'h6073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_143 = 32'h7073 == _control_signal_T_6; // @[Lookup.scala 31:38]
  wire  _control_signal_T_145 = 32'h6b == io_inst; // @[Lookup.scala 31:38]
  wire  _control_signal_T_147 = 32'h7b == io_inst; // @[Lookup.scala 31:38]
  wire  _control_signal_T_148 = _control_signal_T_147 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  wire  _control_signal_T_149 = _control_signal_T_145 ? 1'h0 : _control_signal_T_148; // @[Lookup.scala 33:37]
  wire  _control_signal_T_150 = _control_signal_T_143 ? 1'h0 : _control_signal_T_149; // @[Lookup.scala 33:37]
  wire  _control_signal_T_151 = _control_signal_T_141 ? 1'h0 : _control_signal_T_150; // @[Lookup.scala 33:37]
  wire  _control_signal_T_152 = _control_signal_T_139 ? 1'h0 : _control_signal_T_151; // @[Lookup.scala 33:37]
  wire  _control_signal_T_153 = _control_signal_T_137 ? 1'h0 : _control_signal_T_152; // @[Lookup.scala 33:37]
  wire  _control_signal_T_154 = _control_signal_T_135 ? 1'h0 : _control_signal_T_153; // @[Lookup.scala 33:37]
  wire  _control_signal_T_155 = _control_signal_T_133 ? 1'h0 : _control_signal_T_154; // @[Lookup.scala 33:37]
  wire  _control_signal_T_156 = _control_signal_T_131 ? 1'h0 : _control_signal_T_155; // @[Lookup.scala 33:37]
  wire  _control_signal_T_157 = _control_signal_T_129 ? 1'h0 : _control_signal_T_156; // @[Lookup.scala 33:37]
  wire  _control_signal_T_158 = _control_signal_T_127 ? 1'h0 : _control_signal_T_157; // @[Lookup.scala 33:37]
  wire  _control_signal_T_159 = _control_signal_T_125 ? 1'h0 : _control_signal_T_158; // @[Lookup.scala 33:37]
  wire  _control_signal_T_160 = _control_signal_T_123 ? 1'h0 : _control_signal_T_159; // @[Lookup.scala 33:37]
  wire  _control_signal_T_161 = _control_signal_T_121 ? 1'h0 : _control_signal_T_160; // @[Lookup.scala 33:37]
  wire  _control_signal_T_162 = _control_signal_T_119 ? 1'h0 : _control_signal_T_161; // @[Lookup.scala 33:37]
  wire  _control_signal_T_163 = _control_signal_T_117 ? 1'h0 : _control_signal_T_162; // @[Lookup.scala 33:37]
  wire  _control_signal_T_164 = _control_signal_T_115 ? 1'h0 : _control_signal_T_163; // @[Lookup.scala 33:37]
  wire  _control_signal_T_165 = _control_signal_T_113 ? 1'h0 : _control_signal_T_164; // @[Lookup.scala 33:37]
  wire  _control_signal_T_166 = _control_signal_T_111 ? 1'h0 : _control_signal_T_165; // @[Lookup.scala 33:37]
  wire  _control_signal_T_167 = _control_signal_T_109 ? 1'h0 : _control_signal_T_166; // @[Lookup.scala 33:37]
  wire  _control_signal_T_168 = _control_signal_T_107 ? 1'h0 : _control_signal_T_167; // @[Lookup.scala 33:37]
  wire  _control_signal_T_169 = _control_signal_T_105 ? 1'h0 : _control_signal_T_168; // @[Lookup.scala 33:37]
  wire  _control_signal_T_170 = _control_signal_T_103 ? 1'h0 : _control_signal_T_169; // @[Lookup.scala 33:37]
  wire  _control_signal_T_171 = _control_signal_T_101 ? 1'h0 : _control_signal_T_170; // @[Lookup.scala 33:37]
  wire  _control_signal_T_172 = _control_signal_T_99 ? 1'h0 : _control_signal_T_171; // @[Lookup.scala 33:37]
  wire  _control_signal_T_173 = _control_signal_T_97 ? 1'h0 : _control_signal_T_172; // @[Lookup.scala 33:37]
  wire  _control_signal_T_174 = _control_signal_T_95 ? 1'h0 : _control_signal_T_173; // @[Lookup.scala 33:37]
  wire  _control_signal_T_175 = _control_signal_T_93 ? 1'h0 : _control_signal_T_174; // @[Lookup.scala 33:37]
  wire  _control_signal_T_176 = _control_signal_T_91 ? 1'h0 : _control_signal_T_175; // @[Lookup.scala 33:37]
  wire  _control_signal_T_177 = _control_signal_T_89 ? 1'h0 : _control_signal_T_176; // @[Lookup.scala 33:37]
  wire  _control_signal_T_178 = _control_signal_T_87 ? 1'h0 : _control_signal_T_177; // @[Lookup.scala 33:37]
  wire  _control_signal_T_179 = _control_signal_T_85 ? 1'h0 : _control_signal_T_178; // @[Lookup.scala 33:37]
  wire  _control_signal_T_180 = _control_signal_T_83 ? 1'h0 : _control_signal_T_179; // @[Lookup.scala 33:37]
  wire  _control_signal_T_181 = _control_signal_T_81 ? 1'h0 : _control_signal_T_180; // @[Lookup.scala 33:37]
  wire  _control_signal_T_182 = _control_signal_T_79 ? 1'h0 : _control_signal_T_181; // @[Lookup.scala 33:37]
  wire  _control_signal_T_183 = _control_signal_T_77 ? 1'h0 : _control_signal_T_182; // @[Lookup.scala 33:37]
  wire  _control_signal_T_184 = _control_signal_T_75 ? 1'h0 : _control_signal_T_183; // @[Lookup.scala 33:37]
  wire  _control_signal_T_185 = _control_signal_T_73 ? 1'h0 : _control_signal_T_184; // @[Lookup.scala 33:37]
  wire  _control_signal_T_186 = _control_signal_T_71 ? 1'h0 : _control_signal_T_185; // @[Lookup.scala 33:37]
  wire  _control_signal_T_187 = _control_signal_T_69 ? 1'h0 : _control_signal_T_186; // @[Lookup.scala 33:37]
  wire  _control_signal_T_188 = _control_signal_T_67 ? 1'h0 : _control_signal_T_187; // @[Lookup.scala 33:37]
  wire  _control_signal_T_189 = _control_signal_T_65 ? 1'h0 : _control_signal_T_188; // @[Lookup.scala 33:37]
  wire  _control_signal_T_190 = _control_signal_T_63 ? 1'h0 : _control_signal_T_189; // @[Lookup.scala 33:37]
  wire  _control_signal_T_191 = _control_signal_T_61 ? 1'h0 : _control_signal_T_190; // @[Lookup.scala 33:37]
  wire  _control_signal_T_192 = _control_signal_T_59 ? 1'h0 : _control_signal_T_191; // @[Lookup.scala 33:37]
  wire  _control_signal_T_193 = _control_signal_T_57 ? 1'h0 : _control_signal_T_192; // @[Lookup.scala 33:37]
  wire  _control_signal_T_194 = _control_signal_T_55 ? 1'h0 : _control_signal_T_193; // @[Lookup.scala 33:37]
  wire  _control_signal_T_195 = _control_signal_T_53 ? 1'h0 : _control_signal_T_194; // @[Lookup.scala 33:37]
  wire  _control_signal_T_196 = _control_signal_T_51 ? 1'h0 : _control_signal_T_195; // @[Lookup.scala 33:37]
  wire  _control_signal_T_197 = _control_signal_T_49 ? 1'h0 : _control_signal_T_196; // @[Lookup.scala 33:37]
  wire  _control_signal_T_198 = _control_signal_T_47 ? 1'h0 : _control_signal_T_197; // @[Lookup.scala 33:37]
  wire  _control_signal_T_199 = _control_signal_T_45 ? 1'h0 : _control_signal_T_198; // @[Lookup.scala 33:37]
  wire  _control_signal_T_200 = _control_signal_T_43 ? 1'h0 : _control_signal_T_199; // @[Lookup.scala 33:37]
  wire  _control_signal_T_201 = _control_signal_T_41 ? 1'h0 : _control_signal_T_200; // @[Lookup.scala 33:37]
  wire  _control_signal_T_202 = _control_signal_T_39 ? 1'h0 : _control_signal_T_201; // @[Lookup.scala 33:37]
  wire  _control_signal_T_203 = _control_signal_T_37 ? 1'h0 : _control_signal_T_202; // @[Lookup.scala 33:37]
  wire  _control_signal_T_204 = _control_signal_T_35 ? 1'h0 : _control_signal_T_203; // @[Lookup.scala 33:37]
  wire  _control_signal_T_205 = _control_signal_T_33 ? 1'h0 : _control_signal_T_204; // @[Lookup.scala 33:37]
  wire  _control_signal_T_206 = _control_signal_T_31 ? 1'h0 : _control_signal_T_205; // @[Lookup.scala 33:37]
  wire  _control_signal_T_207 = _control_signal_T_29 ? 1'h0 : _control_signal_T_206; // @[Lookup.scala 33:37]
  wire  _control_signal_T_208 = _control_signal_T_27 ? 1'h0 : _control_signal_T_207; // @[Lookup.scala 33:37]
  wire  _control_signal_T_209 = _control_signal_T_25 ? 1'h0 : _control_signal_T_208; // @[Lookup.scala 33:37]
  wire  _control_signal_T_210 = _control_signal_T_23 ? 1'h0 : _control_signal_T_209; // @[Lookup.scala 33:37]
  wire  _control_signal_T_211 = _control_signal_T_21 ? 1'h0 : _control_signal_T_210; // @[Lookup.scala 33:37]
  wire  _control_signal_T_212 = _control_signal_T_19 ? 1'h0 : _control_signal_T_211; // @[Lookup.scala 33:37]
  wire  _control_signal_T_213 = _control_signal_T_17 ? 1'h0 : _control_signal_T_212; // @[Lookup.scala 33:37]
  wire  _control_signal_T_214 = _control_signal_T_15 ? 1'h0 : _control_signal_T_213; // @[Lookup.scala 33:37]
  wire  _control_signal_T_215 = _control_signal_T_13 ? 1'h0 : _control_signal_T_214; // @[Lookup.scala 33:37]
  wire  _control_signal_T_216 = _control_signal_T_11 ? 1'h0 : _control_signal_T_215; // @[Lookup.scala 33:37]
  wire  _control_signal_T_217 = _control_signal_T_9 ? 1'h0 : _control_signal_T_216; // @[Lookup.scala 33:37]
  wire  _control_signal_T_218 = _control_signal_T_7 ? 1'h0 : _control_signal_T_217; // @[Lookup.scala 33:37]
  wire  _control_signal_T_219 = _control_signal_T_5 ? 1'h0 : _control_signal_T_218; // @[Lookup.scala 33:37]
  wire  _control_signal_T_220 = _control_signal_T_3 ? 1'h0 : _control_signal_T_219; // @[Lookup.scala 33:37]
  wire  control_signal_0 = _control_signal_T_1 ? 1'h0 : _control_signal_T_220; // @[Lookup.scala 33:37]
  wire  _control_signal_T_241 = _control_signal_T_107 | (_control_signal_T_109 | (_control_signal_T_111 | (
    _control_signal_T_113 | (_control_signal_T_115 | (_control_signal_T_117 | (_control_signal_T_119 | (
    _control_signal_T_121 | (_control_signal_T_123 | (_control_signal_T_125 | (_control_signal_T_127 | (
    _control_signal_T_129 | _control_signal_T_131))))))))))); // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_242 = _control_signal_T_105 ? 2'h2 : {{1'd0}, _control_signal_T_241}; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_243 = _control_signal_T_103 ? 2'h2 : _control_signal_T_242; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_244 = _control_signal_T_101 ? 2'h2 : _control_signal_T_243; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_245 = _control_signal_T_99 ? 2'h3 : _control_signal_T_244; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_246 = _control_signal_T_97 ? 2'h3 : _control_signal_T_245; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_247 = _control_signal_T_95 ? 2'h3 : _control_signal_T_246; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_248 = _control_signal_T_93 ? 2'h3 : _control_signal_T_247; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_249 = _control_signal_T_91 ? 2'h3 : _control_signal_T_248; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_250 = _control_signal_T_89 ? 2'h3 : _control_signal_T_249; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_251 = _control_signal_T_87 ? 2'h3 : _control_signal_T_250; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_252 = _control_signal_T_85 ? 2'h3 : _control_signal_T_251; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_253 = _control_signal_T_83 ? 2'h3 : _control_signal_T_252; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_254 = _control_signal_T_81 ? 2'h3 : _control_signal_T_253; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_255 = _control_signal_T_79 ? 2'h3 : _control_signal_T_254; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_256 = _control_signal_T_77 ? 2'h3 : _control_signal_T_255; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_257 = _control_signal_T_75 ? 2'h3 : _control_signal_T_256; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_258 = _control_signal_T_73 ? 2'h3 : _control_signal_T_257; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_259 = _control_signal_T_71 ? 2'h3 : _control_signal_T_258; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_260 = _control_signal_T_69 ? 2'h3 : _control_signal_T_259; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_261 = _control_signal_T_67 ? 2'h3 : _control_signal_T_260; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_262 = _control_signal_T_65 ? 2'h3 : _control_signal_T_261; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_263 = _control_signal_T_63 ? 2'h3 : _control_signal_T_262; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_264 = _control_signal_T_61 ? 2'h3 : _control_signal_T_263; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_265 = _control_signal_T_59 ? 2'h3 : _control_signal_T_264; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_266 = _control_signal_T_57 ? 2'h3 : _control_signal_T_265; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_267 = _control_signal_T_55 ? 2'h0 : _control_signal_T_266; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_268 = _control_signal_T_53 ? 2'h0 : _control_signal_T_267; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_269 = _control_signal_T_51 ? 2'h0 : _control_signal_T_268; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_270 = _control_signal_T_49 ? 2'h3 : _control_signal_T_269; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_271 = _control_signal_T_47 ? 2'h3 : _control_signal_T_270; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_272 = _control_signal_T_45 ? 2'h3 : _control_signal_T_271; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_273 = _control_signal_T_43 ? 2'h3 : _control_signal_T_272; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_274 = _control_signal_T_41 ? 2'h3 : _control_signal_T_273; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_275 = _control_signal_T_39 ? 2'h3 : _control_signal_T_274; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_276 = _control_signal_T_37 ? 2'h2 : _control_signal_T_275; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_277 = _control_signal_T_35 ? 2'h2 : _control_signal_T_276; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_278 = _control_signal_T_33 ? 2'h2 : _control_signal_T_277; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_279 = _control_signal_T_31 ? 2'h2 : _control_signal_T_278; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_280 = _control_signal_T_29 ? 2'h2 : _control_signal_T_279; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_281 = _control_signal_T_27 ? 2'h2 : _control_signal_T_280; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_282 = _control_signal_T_25 ? 2'h2 : _control_signal_T_281; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_283 = _control_signal_T_23 ? 2'h2 : _control_signal_T_282; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_284 = _control_signal_T_21 ? 2'h0 : _control_signal_T_283; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_285 = _control_signal_T_19 ? 2'h0 : _control_signal_T_284; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_286 = _control_signal_T_17 ? 2'h0 : _control_signal_T_285; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_287 = _control_signal_T_15 ? 2'h0 : _control_signal_T_286; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_288 = _control_signal_T_13 ? 2'h0 : _control_signal_T_287; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_289 = _control_signal_T_11 ? 2'h0 : _control_signal_T_288; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_290 = _control_signal_T_9 ? 2'h0 : _control_signal_T_289; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_291 = _control_signal_T_7 ? 2'h0 : _control_signal_T_290; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_292 = _control_signal_T_5 ? 2'h0 : _control_signal_T_291; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_293 = _control_signal_T_3 ? 2'h3 : _control_signal_T_292; // @[Lookup.scala 33:37]
  wire [1:0] control_signal_1 = _control_signal_T_1 ? 2'h3 : _control_signal_T_293; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_85 = _control_signal_T_3 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] alu_signal_0 = _control_signal_T_1 ? 2'h0 : _alu_signal_T_85; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_91 = _control_signal_T_89 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_92 = _control_signal_T_87 ? 2'h1 : _alu_signal_T_91; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_93 = _control_signal_T_85 ? 2'h1 : _alu_signal_T_92; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_94 = _control_signal_T_83 ? 2'h1 : _alu_signal_T_93; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_95 = _control_signal_T_81 ? 2'h1 : _alu_signal_T_94; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_96 = _control_signal_T_79 ? 2'h1 : _alu_signal_T_95; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_97 = _control_signal_T_77 ? 2'h1 : _alu_signal_T_96; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_98 = _control_signal_T_49 ? 2'h1 : _alu_signal_T_97; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_99 = _control_signal_T_47 ? 2'h1 : _alu_signal_T_98; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_100 = _control_signal_T_45 ? 2'h1 : _alu_signal_T_99; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_101 = _control_signal_T_43 ? 2'h1 : _alu_signal_T_100; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_102 = _control_signal_T_41 ? 2'h1 : _alu_signal_T_101; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_103 = _control_signal_T_39 ? 2'h1 : _alu_signal_T_102; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_104 = _control_signal_T_75 ? 2'h0 : _alu_signal_T_103; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_105 = _control_signal_T_73 ? 2'h0 : _alu_signal_T_104; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_106 = _control_signal_T_71 ? 2'h0 : _alu_signal_T_105; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_107 = _control_signal_T_69 ? 2'h0 : _alu_signal_T_106; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_108 = _control_signal_T_67 ? 2'h0 : _alu_signal_T_107; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_109 = _control_signal_T_65 ? 2'h0 : _alu_signal_T_108; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_110 = _control_signal_T_63 ? 2'h0 : _alu_signal_T_109; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_111 = _control_signal_T_61 ? 2'h0 : _alu_signal_T_110; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_112 = _control_signal_T_59 ? 2'h0 : _alu_signal_T_111; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_113 = _control_signal_T_3 ? 2'h1 : _alu_signal_T_112; // @[Lookup.scala 33:37]
  wire [1:0] alu_signal_1 = _control_signal_T_1 ? 2'h1 : _alu_signal_T_113; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_114 = _control_signal_T_99 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_115 = _control_signal_T_97 ? 4'h8 : _alu_signal_T_114; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_116 = _control_signal_T_95 ? 4'h7 : _alu_signal_T_115; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_117 = _control_signal_T_93 ? 4'h1 : _alu_signal_T_116; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_118 = _control_signal_T_91 ? 4'h0 : _alu_signal_T_117; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_119 = _control_signal_T_89 ? 4'h9 : _alu_signal_T_118; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_120 = _control_signal_T_87 ? 4'h8 : _alu_signal_T_119; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_121 = _control_signal_T_85 ? 4'h7 : _alu_signal_T_120; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_122 = _control_signal_T_83 ? 4'h0 : _alu_signal_T_121; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_123 = _control_signal_T_81 ? 4'h9 : _alu_signal_T_122; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_124 = _control_signal_T_79 ? 4'h8 : _alu_signal_T_123; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_125 = _control_signal_T_77 ? 4'h7 : _alu_signal_T_124; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_126 = _control_signal_T_49 ? 4'h5 : _alu_signal_T_125; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_127 = _control_signal_T_47 ? 4'h6 : _alu_signal_T_126; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_128 = _control_signal_T_45 ? 4'h4 : _alu_signal_T_127; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_129 = _control_signal_T_43 ? 4'h3 : _alu_signal_T_128; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_130 = _control_signal_T_41 ? 4'h2 : _alu_signal_T_129; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_131 = _control_signal_T_39 ? 4'h0 : _alu_signal_T_130; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_132 = _control_signal_T_75 ? 4'h5 : _alu_signal_T_131; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_133 = _control_signal_T_73 ? 4'h6 : _alu_signal_T_132; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_134 = _control_signal_T_71 ? 4'h9 : _alu_signal_T_133; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_135 = _control_signal_T_69 ? 4'h8 : _alu_signal_T_134; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_136 = _control_signal_T_67 ? 4'h4 : _alu_signal_T_135; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_137 = _control_signal_T_65 ? 4'h3 : _alu_signal_T_136; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_138 = _control_signal_T_63 ? 4'h2 : _alu_signal_T_137; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_139 = _control_signal_T_61 ? 4'h7 : _alu_signal_T_138; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_140 = _control_signal_T_59 ? 4'h1 : _alu_signal_T_139; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_141 = _control_signal_T_3 ? 4'h0 : _alu_signal_T_140; // @[Lookup.scala 33:37]
  wire [3:0] alu_signal_2 = _control_signal_T_1 ? 4'ha : _alu_signal_T_141; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_147 = _control_signal_T_89 ? shamtIMM : 20'h0; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_148 = _control_signal_T_87 ? shamtIMM : _alu_signal_T_147; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_149 = _control_signal_T_85 ? shamtIMM : _alu_signal_T_148; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_150 = _control_signal_T_83 ? aluIIMM : _alu_signal_T_149; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_151 = _control_signal_T_81 ? shamtIMM : _alu_signal_T_150; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_152 = _control_signal_T_79 ? shamtIMM : _alu_signal_T_151; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_153 = _control_signal_T_77 ? shamtIMM : _alu_signal_T_152; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_154 = _control_signal_T_49 ? aluIIMM : _alu_signal_T_153; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_155 = _control_signal_T_47 ? aluIIMM : _alu_signal_T_154; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_156 = _control_signal_T_45 ? aluIIMM : _alu_signal_T_155; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_157 = _control_signal_T_43 ? aluIIMM : _alu_signal_T_156; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_158 = _control_signal_T_41 ? aluIIMM : _alu_signal_T_157; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_159 = _control_signal_T_39 ? aluIIMM : _alu_signal_T_158; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_160 = _control_signal_T_75 ? 20'h0 : _alu_signal_T_159; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_161 = _control_signal_T_73 ? 20'h0 : _alu_signal_T_160; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_162 = _control_signal_T_71 ? 20'h0 : _alu_signal_T_161; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_163 = _control_signal_T_69 ? 20'h0 : _alu_signal_T_162; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_164 = _control_signal_T_67 ? 20'h0 : _alu_signal_T_163; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_165 = _control_signal_T_65 ? 20'h0 : _alu_signal_T_164; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_166 = _control_signal_T_63 ? 20'h0 : _alu_signal_T_165; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_167 = _control_signal_T_61 ? 20'h0 : _alu_signal_T_166; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_168 = _control_signal_T_59 ? 20'h0 : _alu_signal_T_167; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_169 = _control_signal_T_3 ? aluUIMM : _alu_signal_T_168; // @[Lookup.scala 33:37]
  wire [19:0] alu_signal_3 = _control_signal_T_1 ? aluUIMM : _alu_signal_T_169; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_179 = _control_signal_T_81 ? 1'h0 : _control_signal_T_83 | (_control_signal_T_85 | (
    _control_signal_T_87 | (_control_signal_T_89 | (_control_signal_T_91 | (_control_signal_T_93 | (_control_signal_T_95
     | (_control_signal_T_97 | _control_signal_T_99))))))); // @[Lookup.scala 33:37]
  wire  _alu_signal_T_180 = _control_signal_T_79 ? 1'h0 : _alu_signal_T_179; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_181 = _control_signal_T_77 ? 1'h0 : _alu_signal_T_180; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_182 = _control_signal_T_49 ? 1'h0 : _alu_signal_T_181; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_183 = _control_signal_T_47 ? 1'h0 : _alu_signal_T_182; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_184 = _control_signal_T_45 ? 1'h0 : _alu_signal_T_183; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_185 = _control_signal_T_43 ? 1'h0 : _alu_signal_T_184; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_186 = _control_signal_T_41 ? 1'h0 : _alu_signal_T_185; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_187 = _control_signal_T_39 ? 1'h0 : _alu_signal_T_186; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_188 = _control_signal_T_75 ? 1'h0 : _alu_signal_T_187; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_189 = _control_signal_T_73 ? 1'h0 : _alu_signal_T_188; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_190 = _control_signal_T_71 ? 1'h0 : _alu_signal_T_189; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_191 = _control_signal_T_69 ? 1'h0 : _alu_signal_T_190; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_192 = _control_signal_T_67 ? 1'h0 : _alu_signal_T_191; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_193 = _control_signal_T_65 ? 1'h0 : _alu_signal_T_192; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_194 = _control_signal_T_63 ? 1'h0 : _alu_signal_T_193; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_195 = _control_signal_T_61 ? 1'h0 : _alu_signal_T_194; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_196 = _control_signal_T_59 ? 1'h0 : _alu_signal_T_195; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_197 = _control_signal_T_3 ? 1'h0 : _alu_signal_T_196; // @[Lookup.scala 33:37]
  wire  alu_signal_4 = _control_signal_T_1 ? 1'h0 : _alu_signal_T_197; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_225 = _control_signal_T_3 ? 5'h0 : IRS; // @[Lookup.scala 33:37]
  wire [4:0] alu_signal_5 = _control_signal_T_1 ? 5'h0 : _alu_signal_T_225; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_231 = _control_signal_T_89 ? 5'h0 : IRT; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_232 = _control_signal_T_87 ? 5'h0 : _alu_signal_T_231; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_233 = _control_signal_T_85 ? 5'h0 : _alu_signal_T_232; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_234 = _control_signal_T_83 ? 5'h0 : _alu_signal_T_233; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_235 = _control_signal_T_81 ? 5'h0 : _alu_signal_T_234; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_236 = _control_signal_T_79 ? 5'h0 : _alu_signal_T_235; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_237 = _control_signal_T_77 ? 5'h0 : _alu_signal_T_236; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_238 = _control_signal_T_49 ? 5'h0 : _alu_signal_T_237; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_239 = _control_signal_T_47 ? 5'h0 : _alu_signal_T_238; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_240 = _control_signal_T_45 ? 5'h0 : _alu_signal_T_239; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_241 = _control_signal_T_43 ? 5'h0 : _alu_signal_T_240; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_242 = _control_signal_T_41 ? 5'h0 : _alu_signal_T_241; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_243 = _control_signal_T_39 ? 5'h0 : _alu_signal_T_242; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_244 = _control_signal_T_75 ? IRT : _alu_signal_T_243; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_245 = _control_signal_T_73 ? IRT : _alu_signal_T_244; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_246 = _control_signal_T_71 ? IRT : _alu_signal_T_245; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_247 = _control_signal_T_69 ? IRT : _alu_signal_T_246; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_248 = _control_signal_T_67 ? IRT : _alu_signal_T_247; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_249 = _control_signal_T_65 ? IRT : _alu_signal_T_248; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_250 = _control_signal_T_63 ? IRT : _alu_signal_T_249; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_251 = _control_signal_T_61 ? IRT : _alu_signal_T_250; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_252 = _control_signal_T_59 ? IRT : _alu_signal_T_251; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_253 = _control_signal_T_3 ? 5'h0 : _alu_signal_T_252; // @[Lookup.scala 33:37]
  wire [4:0] alu_signal_6 = _control_signal_T_1 ? 5'h0 : _alu_signal_T_253; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_24 = _control_signal_T_131 ? 5'h17 : 5'h14; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_25 = _control_signal_T_129 ? 5'h16 : _mdu_signal_T_24; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_26 = _control_signal_T_127 ? 5'h15 : _mdu_signal_T_25; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_27 = _control_signal_T_125 ? 5'h14 : _mdu_signal_T_26; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_28 = _control_signal_T_123 ? 5'h10 : _mdu_signal_T_27; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_29 = _control_signal_T_121 ? 5'h17 : _mdu_signal_T_28; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_30 = _control_signal_T_119 ? 5'h16 : _mdu_signal_T_29; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_31 = _control_signal_T_117 ? 5'h15 : _mdu_signal_T_30; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_32 = _control_signal_T_113 ? 5'h12 : _mdu_signal_T_31; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_33 = _control_signal_T_111 ? 5'h13 : _mdu_signal_T_32; // @[Lookup.scala 33:37]
  wire [4:0] _mdu_signal_T_34 = _control_signal_T_109 ? 5'h11 : _mdu_signal_T_33; // @[Lookup.scala 33:37]
  wire [4:0] mdu_signal_0 = _control_signal_T_107 ? 5'h10 : _mdu_signal_T_34; // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_40 = _control_signal_T_121 ? 1'h0 : _control_signal_T_123 | (_control_signal_T_125 | (
    _control_signal_T_127 | (_control_signal_T_129 | _control_signal_T_131))); // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_41 = _control_signal_T_119 ? 1'h0 : _mdu_signal_T_40; // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_42 = _control_signal_T_117 ? 1'h0 : _mdu_signal_T_41; // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_43 = _control_signal_T_113 ? 1'h0 : _mdu_signal_T_42; // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_44 = _control_signal_T_111 ? 1'h0 : _mdu_signal_T_43; // @[Lookup.scala 33:37]
  wire  _mdu_signal_T_45 = _control_signal_T_109 ? 1'h0 : _mdu_signal_T_44; // @[Lookup.scala 33:37]
  wire  mdu_signal_1 = _control_signal_T_107 ? 1'h0 : _mdu_signal_T_45; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_21 = _control_signal_T_105 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_23 = _control_signal_T_37 ? 1'h0 : _control_signal_T_101 | _lsu_signal_T_21; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_24 = _control_signal_T_35 ? 1'h0 : _lsu_signal_T_23; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_25 = _control_signal_T_33 ? 1'h0 : _lsu_signal_T_24; // @[Lookup.scala 33:37]
  wire  lsu_signal_0 = _control_signal_T_25 | (_control_signal_T_27 | (_control_signal_T_29 | (_control_signal_T_31 |
    _lsu_signal_T_25))); // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_29 = _control_signal_T_103 ? 3'h6 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_30 = _control_signal_T_105 ? 3'h5 : _lsu_signal_T_29; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_31 = _control_signal_T_101 ? 3'h5 : _lsu_signal_T_30; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_32 = _control_signal_T_37 ? 3'h4 : _lsu_signal_T_31; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_33 = _control_signal_T_35 ? 3'h2 : _lsu_signal_T_32; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_34 = _control_signal_T_33 ? 3'h0 : _lsu_signal_T_33; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_35 = _control_signal_T_31 ? 3'h3 : _lsu_signal_T_34; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_36 = _control_signal_T_29 ? 3'h1 : _lsu_signal_T_35; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_37 = _control_signal_T_27 ? 3'h4 : _lsu_signal_T_36; // @[Lookup.scala 33:37]
  wire [2:0] lsu_signal_1 = _control_signal_T_25 ? 3'h2 : _lsu_signal_T_37; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_39 = _control_signal_T_105 ? 5'h0 : IRD; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_40 = _control_signal_T_101 ? IRD : _lsu_signal_T_39; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_41 = _control_signal_T_37 ? 5'h0 : _lsu_signal_T_40; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_42 = _control_signal_T_35 ? 5'h0 : _lsu_signal_T_41; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_43 = _control_signal_T_33 ? 5'h0 : _lsu_signal_T_42; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_44 = _control_signal_T_31 ? IRD : _lsu_signal_T_43; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_45 = _control_signal_T_29 ? IRD : _lsu_signal_T_44; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_46 = _control_signal_T_27 ? IRD : _lsu_signal_T_45; // @[Lookup.scala 33:37]
  wire [4:0] lsu_signal_2 = _control_signal_T_25 ? IRD : _lsu_signal_T_46; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_57 = _control_signal_T_105 ? IRT : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_58 = _control_signal_T_101 ? 5'h0 : _lsu_signal_T_57; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_59 = _control_signal_T_37 ? IRT : _lsu_signal_T_58; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_60 = _control_signal_T_35 ? IRT : _lsu_signal_T_59; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_61 = _control_signal_T_33 ? IRT : _lsu_signal_T_60; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_62 = _control_signal_T_31 ? 5'h0 : _lsu_signal_T_61; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_63 = _control_signal_T_29 ? 5'h0 : _lsu_signal_T_62; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_64 = _control_signal_T_27 ? 5'h0 : _lsu_signal_T_63; // @[Lookup.scala 33:37]
  wire [4:0] lsu_signal_4 = _control_signal_T_25 ? 5'h0 : _lsu_signal_T_64; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_38 = _control_signal_T_147 ? 4'h3 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_39 = _control_signal_T_145 ? 4'h3 : _bju_signal_T_38; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_40 = _control_signal_T_143 ? 4'h0 : _bju_signal_T_39; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_41 = _control_signal_T_141 ? 4'h0 : _bju_signal_T_40; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_42 = _control_signal_T_139 ? 4'h0 : _bju_signal_T_41; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_43 = _control_signal_T_137 ? 4'h0 : _bju_signal_T_42; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_44 = _control_signal_T_135 ? 4'h0 : _bju_signal_T_43; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_45 = _control_signal_T_133 ? 4'h0 : _bju_signal_T_44; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_46 = _control_signal_T_53 ? 4'h7 : _bju_signal_T_45; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_47 = _control_signal_T_51 ? 4'h6 : _bju_signal_T_46; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_48 = _control_signal_T_21 ? 4'h5 : _bju_signal_T_47; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_49 = _control_signal_T_7 ? 4'h4 : _bju_signal_T_48; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_50 = _control_signal_T_5 ? 4'h3 : _bju_signal_T_49; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_51 = _control_signal_T_19 ? 4'h2 : _bju_signal_T_50; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_52 = _control_signal_T_17 ? 4'h2 : _bju_signal_T_51; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_53 = _control_signal_T_15 ? 4'h2 : _bju_signal_T_52; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_54 = _control_signal_T_13 ? 4'h2 : _bju_signal_T_53; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_55 = _control_signal_T_11 ? 4'h2 : _bju_signal_T_54; // @[Lookup.scala 33:37]
  wire [3:0] bju_signal_0 = _control_signal_T_9 ? 4'h2 : _bju_signal_T_55; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_58 = _control_signal_T_143 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_59 = _control_signal_T_141 ? 2'h1 : _bju_signal_T_58; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_60 = _control_signal_T_139 ? 2'h1 : _bju_signal_T_59; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_61 = _control_signal_T_137 ? 2'h0 : _bju_signal_T_60; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_62 = _control_signal_T_135 ? 2'h0 : _bju_signal_T_61; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_63 = _control_signal_T_133 ? 2'h0 : _bju_signal_T_62; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_64 = _control_signal_T_53 ? 2'h0 : _bju_signal_T_63; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_65 = _control_signal_T_51 ? 2'h0 : _bju_signal_T_64; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_66 = _control_signal_T_21 ? 2'h0 : _bju_signal_T_65; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_67 = _control_signal_T_7 ? 2'h0 : _bju_signal_T_66; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_68 = _control_signal_T_5 ? 2'h0 : _bju_signal_T_67; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_69 = _control_signal_T_19 ? 2'h0 : _bju_signal_T_68; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_70 = _control_signal_T_17 ? 2'h0 : _bju_signal_T_69; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_71 = _control_signal_T_15 ? 2'h0 : _bju_signal_T_70; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_72 = _control_signal_T_13 ? 2'h0 : _bju_signal_T_71; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_73 = _control_signal_T_11 ? 2'h0 : _bju_signal_T_72; // @[Lookup.scala 33:37]
  wire [1:0] bju_signal_1 = _control_signal_T_9 ? 2'h0 : _bju_signal_T_73; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_74 = _control_signal_T_147 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_75 = _control_signal_T_145 ? 2'h1 : _bju_signal_T_74; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_76 = _control_signal_T_143 ? 2'h2 : _bju_signal_T_75; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_77 = _control_signal_T_141 ? 2'h2 : _bju_signal_T_76; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_78 = _control_signal_T_139 ? 2'h2 : _bju_signal_T_77; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_79 = _control_signal_T_137 ? 2'h2 : _bju_signal_T_78; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_80 = _control_signal_T_135 ? 2'h2 : _bju_signal_T_79; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_81 = _control_signal_T_133 ? 2'h2 : _bju_signal_T_80; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_82 = _control_signal_T_53 ? 2'h0 : _bju_signal_T_81; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_83 = _control_signal_T_51 ? 2'h0 : _bju_signal_T_82; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_84 = _control_signal_T_21 ? 2'h0 : _bju_signal_T_83; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_85 = _control_signal_T_7 ? 2'h1 : _bju_signal_T_84; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_86 = _control_signal_T_5 ? 2'h1 : _bju_signal_T_85; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_87 = _control_signal_T_19 ? 2'h0 : _bju_signal_T_86; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_88 = _control_signal_T_17 ? 2'h0 : _bju_signal_T_87; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_89 = _control_signal_T_15 ? 2'h0 : _bju_signal_T_88; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_90 = _control_signal_T_13 ? 2'h0 : _bju_signal_T_89; // @[Lookup.scala 33:37]
  wire [1:0] _bju_signal_T_91 = _control_signal_T_11 ? 2'h0 : _bju_signal_T_90; // @[Lookup.scala 33:37]
  wire [1:0] bju_signal_2 = _control_signal_T_9 ? 2'h0 : _bju_signal_T_91; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_100 = _control_signal_T_53 ? 1'h0 : _control_signal_T_133 | (_control_signal_T_135 | (
    _control_signal_T_137 | (_control_signal_T_139 | (_control_signal_T_141 | (_control_signal_T_143 | (
    _control_signal_T_145 | _control_signal_T_147)))))); // @[Lookup.scala 33:37]
  wire  _bju_signal_T_101 = _control_signal_T_51 ? 1'h0 : _bju_signal_T_100; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_102 = _control_signal_T_21 ? 1'h0 : _bju_signal_T_101; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_105 = _control_signal_T_19 ? 1'h0 : _control_signal_T_5 | (_control_signal_T_7 | _bju_signal_T_102
    ); // @[Lookup.scala 33:37]
  wire  _bju_signal_T_106 = _control_signal_T_17 ? 1'h0 : _bju_signal_T_105; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_107 = _control_signal_T_15 ? 1'h0 : _bju_signal_T_106; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_108 = _control_signal_T_13 ? 1'h0 : _bju_signal_T_107; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_109 = _control_signal_T_11 ? 1'h0 : _bju_signal_T_108; // @[Lookup.scala 33:37]
  wire  bju_signal_3 = _control_signal_T_9 ? 1'h0 : _bju_signal_T_109; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_112 = _control_signal_T_143 ? 4'hb : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_113 = _control_signal_T_141 ? 4'h6 : _bju_signal_T_112; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_114 = _control_signal_T_139 ? 4'h0 : _bju_signal_T_113; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_115 = _control_signal_T_137 ? 4'hb : _bju_signal_T_114; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_116 = _control_signal_T_135 ? 4'h6 : _bju_signal_T_115; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_117 = _control_signal_T_133 ? 4'h0 : _bju_signal_T_116; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_118 = _control_signal_T_53 ? 4'h0 : _bju_signal_T_117; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_119 = _control_signal_T_51 ? 4'h0 : _bju_signal_T_118; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_120 = _control_signal_T_21 ? 4'h0 : _bju_signal_T_119; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_121 = _control_signal_T_7 ? 4'h0 : _bju_signal_T_120; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_122 = _control_signal_T_5 ? 4'h0 : _bju_signal_T_121; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_123 = _control_signal_T_19 ? 4'h3 : _bju_signal_T_122; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_124 = _control_signal_T_17 ? 4'h3 : _bju_signal_T_123; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_125 = _control_signal_T_15 ? 4'h1 : _bju_signal_T_124; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_126 = _control_signal_T_13 ? 4'h1 : _bju_signal_T_125; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_127 = _control_signal_T_11 ? 4'h1 : _bju_signal_T_126; // @[Lookup.scala 33:37]
  wire [3:0] bju_signal_4 = _control_signal_T_9 ? 4'h1 : _bju_signal_T_127; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_128 = _control_signal_T_147 ? 64'h4 : 64'h0; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_129 = _control_signal_T_145 ? 64'h0 : _bju_signal_T_128; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_130 = _control_signal_T_143 ? {{44'd0}, CSRIMM} : _bju_signal_T_129; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_131 = _control_signal_T_141 ? {{44'd0}, CSRIMM} : _bju_signal_T_130; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_132 = _control_signal_T_139 ? {{44'd0}, CSRIMM} : _bju_signal_T_131; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_133 = _control_signal_T_137 ? {{44'd0}, CSRIMM} : _bju_signal_T_132; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_134 = _control_signal_T_135 ? {{44'd0}, CSRIMM} : _bju_signal_T_133; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_135 = _control_signal_T_133 ? {{44'd0}, CSRIMM} : _bju_signal_T_134; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_136 = _control_signal_T_53 ? 64'h0 : _bju_signal_T_135; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_137 = _control_signal_T_51 ? 64'h0 : _bju_signal_T_136; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_138 = _control_signal_T_21 ? 64'h0 : _bju_signal_T_137; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_139 = _control_signal_T_7 ? {{44'd0}, aluIIMM} : _bju_signal_T_138; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_140 = _control_signal_T_5 ? {{44'd0}, JIMM} : _bju_signal_T_139; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_141 = _control_signal_T_19 ? {{44'd0}, BIMM} : _bju_signal_T_140; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_142 = _control_signal_T_17 ? {{44'd0}, BIMM} : _bju_signal_T_141; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_143 = _control_signal_T_15 ? {{44'd0}, BIMM} : _bju_signal_T_142; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_144 = _control_signal_T_13 ? {{44'd0}, BIMM} : _bju_signal_T_143; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_145 = _control_signal_T_11 ? {{44'd0}, BIMM} : _bju_signal_T_144; // @[Lookup.scala 33:37]
  wire [63:0] bju_signal_5 = _control_signal_T_9 ? {{44'd0}, BIMM} : _bju_signal_T_145; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_148 = _control_signal_T_143 ? IRD : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_149 = _control_signal_T_141 ? IRD : _bju_signal_T_148; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_150 = _control_signal_T_139 ? IRD : _bju_signal_T_149; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_151 = _control_signal_T_137 ? IRD : _bju_signal_T_150; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_152 = _control_signal_T_135 ? IRD : _bju_signal_T_151; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_153 = _control_signal_T_133 ? IRD : _bju_signal_T_152; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_154 = _control_signal_T_53 ? 5'h0 : _bju_signal_T_153; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_155 = _control_signal_T_51 ? 5'h0 : _bju_signal_T_154; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_156 = _control_signal_T_21 ? 5'h0 : _bju_signal_T_155; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_157 = _control_signal_T_7 ? IRD : _bju_signal_T_156; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_158 = _control_signal_T_5 ? IRD : _bju_signal_T_157; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_159 = _control_signal_T_19 ? 5'h0 : _bju_signal_T_158; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_160 = _control_signal_T_17 ? 5'h0 : _bju_signal_T_159; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_161 = _control_signal_T_15 ? 5'h0 : _bju_signal_T_160; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_162 = _control_signal_T_13 ? 5'h0 : _bju_signal_T_161; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_163 = _control_signal_T_11 ? 5'h0 : _bju_signal_T_162; // @[Lookup.scala 33:37]
  wire [4:0] bju_signal_6 = _control_signal_T_9 ? 5'h0 : _bju_signal_T_163; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_166 = _control_signal_T_143 ? IRS : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_167 = _control_signal_T_141 ? IRS : _bju_signal_T_166; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_168 = _control_signal_T_139 ? IRS : _bju_signal_T_167; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_169 = _control_signal_T_137 ? IRS : _bju_signal_T_168; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_170 = _control_signal_T_135 ? IRS : _bju_signal_T_169; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_171 = _control_signal_T_133 ? IRS : _bju_signal_T_170; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_172 = _control_signal_T_53 ? 5'h0 : _bju_signal_T_171; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_173 = _control_signal_T_51 ? 5'h0 : _bju_signal_T_172; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_174 = _control_signal_T_21 ? 5'h0 : _bju_signal_T_173; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_175 = _control_signal_T_7 ? IRS : _bju_signal_T_174; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_176 = _control_signal_T_5 ? 5'h0 : _bju_signal_T_175; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_177 = _control_signal_T_19 ? IRS : _bju_signal_T_176; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_178 = _control_signal_T_17 ? IRS : _bju_signal_T_177; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_179 = _control_signal_T_15 ? IRS : _bju_signal_T_178; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_180 = _control_signal_T_13 ? IRS : _bju_signal_T_179; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_181 = _control_signal_T_11 ? IRS : _bju_signal_T_180; // @[Lookup.scala 33:37]
  wire [4:0] bju_signal_7 = _control_signal_T_9 ? IRS : _bju_signal_T_181; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_195 = _control_signal_T_19 ? IRT : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_196 = _control_signal_T_17 ? IRT : _bju_signal_T_195; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_197 = _control_signal_T_15 ? IRT : _bju_signal_T_196; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_198 = _control_signal_T_13 ? IRT : _bju_signal_T_197; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_199 = _control_signal_T_11 ? IRT : _bju_signal_T_198; // @[Lookup.scala 33:37]
  wire [4:0] bju_signal_8 = _control_signal_T_9 ? IRT : _bju_signal_T_199; // @[Lookup.scala 33:37]
  wire [3:0] _branch_signal_T_12 = _control_signal_T_19 ? 4'h5 : 4'h1; // @[Lookup.scala 33:37]
  wire [3:0] _branch_signal_T_13 = _control_signal_T_17 ? 4'h4 : _branch_signal_T_12; // @[Lookup.scala 33:37]
  wire [3:0] _branch_signal_T_14 = _control_signal_T_15 ? 4'h3 : _branch_signal_T_13; // @[Lookup.scala 33:37]
  wire [3:0] _branch_signal_T_15 = _control_signal_T_13 ? 4'h6 : _branch_signal_T_14; // @[Lookup.scala 33:37]
  wire [3:0] _branch_signal_T_16 = _control_signal_T_11 ? 4'h2 : _branch_signal_T_15; // @[Lookup.scala 33:37]
  wire [3:0] branch_signal_0 = _control_signal_T_9 ? 4'h1 : _branch_signal_T_16; // @[Lookup.scala 33:37]
  wire  _io_mops_branch_type_T = control_signal_1 == 2'h0; // @[Decode.scala 314:50]
  wire [1:0] _io_mops_src_a_T_1 = 2'h3 == control_signal_1 ? alu_signal_0 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] _io_mops_src_b_T_1 = 2'h3 == control_signal_1 ? alu_signal_1 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] _io_mops_src_b_T_3 = 2'h0 == control_signal_1 ? bju_signal_2 : _io_mops_src_b_T_1; // @[Mux.scala 80:57]
  wire  _io_mops_write_dest_T_1 = 2'h2 == control_signal_1 ? lsu_signal_0 : 1'h1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_alu_op_T_1 = 2'h1 == control_signal_1 ? mdu_signal_0 : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_alu_op_T_3 = 2'h3 == control_signal_1 ? {{1'd0}, alu_signal_2} : _io_mops_alu_op_T_1; // @[Mux.scala 80:57]
  wire [1:0] _io_mops_write_src_T_3 = bju_signal_0 == 4'h3 | bju_signal_0 == 4'h4 ? 2'h3 : 2'h0; // @[Decode.scala 352:21]
  wire [1:0] _io_mops_write_src_T_5 = 2'h2 == control_signal_1 ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs1_T_1 = 2'h1 == control_signal_1 ? IRS : alu_signal_5; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs1_T_3 = 2'h0 == control_signal_1 ? bju_signal_7 : _io_mops_rs1_T_1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs2_T_1 = 2'h1 == control_signal_1 ? IRT : alu_signal_6; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs2_T_3 = 2'h0 == control_signal_1 ? bju_signal_8 : _io_mops_rs2_T_1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rd_T_3 = 2'h0 == control_signal_1 ? bju_signal_6 : IRD; // @[Mux.scala 80:57]
  wire [19:0] _io_mops_imm_T_1 = ~lsu_signal_0 ? lsuSIMM : aluIIMM; // @[Mux.scala 80:57]
  wire [19:0] _io_mops_imm_T_3 = 2'h3 == control_signal_1 ? alu_signal_3 : _io_mops_imm_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_mops_imm_T_5 = 2'h0 == control_signal_1 ? bju_signal_5 : {{44'd0}, _io_mops_imm_T_3}; // @[Mux.scala 80:57]
  assign io_mops_illegal = control_signal_0 | |io_pc[1:0]; // @[Decode.scala 313:53]
  assign io_mops_next_pc = _io_mops_branch_type_T ? bju_signal_0 : 4'h0; // @[Decode.scala 316:31]
  assign io_mops_alu_mdu_lsu = _control_signal_T_1 ? 2'h3 : _control_signal_T_293; // @[Lookup.scala 33:37]
  assign io_mops_branch_type = control_signal_1 == 2'h0 & bju_signal_0 == 4'h2 ? branch_signal_0 : 4'h0; // @[Decode.scala 314:31]
  assign io_mops_src_a = 2'h0 == control_signal_1 ? bju_signal_1 : _io_mops_src_a_T_1; // @[Mux.scala 80:57]
  assign io_mops_src_b = 2'h2 == control_signal_1 ? 2'h1 : _io_mops_src_b_T_3; // @[Mux.scala 80:57]
  assign io_mops_write_dest = 2'h0 == control_signal_1 ? bju_signal_3 : _io_mops_write_dest_T_1; // @[Mux.scala 80:57]
  assign io_mops_alu_op = 2'h0 == control_signal_1 ? {{1'd0}, bju_signal_4} : _io_mops_alu_op_T_3; // @[Mux.scala 80:57]
  assign io_mops_alu_expand = 2'h1 == control_signal_1 ? mdu_signal_1 : alu_signal_4; // @[Mux.scala 80:57]
  assign io_mops_mem_width = control_signal_1 == 2'h2 ? lsu_signal_1 : 3'h0; // @[Decode.scala 348:31]
  assign io_mops_write_src = 2'h0 == control_signal_1 ? _io_mops_write_src_T_3 : _io_mops_write_src_T_5; // @[Mux.scala 80:57]
  assign io_mops_rs1 = 2'h2 == control_signal_1 ? IRS : _io_mops_rs1_T_3; // @[Mux.scala 80:57]
  assign io_mops_rs2 = 2'h2 == control_signal_1 ? lsu_signal_4 : _io_mops_rs2_T_3; // @[Mux.scala 80:57]
  assign io_mops_rd = 2'h2 == control_signal_1 ? lsu_signal_2 : _io_mops_rd_T_3; // @[Mux.scala 80:57]
  assign io_mops_imm = _io_mops_imm_T_5[19:0]; // @[Decode.scala 376:25]
  assign io_mops_pc = io_pc; // @[Decode.scala 383:25]
  assign io_mops_predict_taken = io_bht_predict_taken; // @[Decode.scala 384:25]
  assign io_mops_target_pc = io_target_pc; // @[Decode.scala 385:25]
  assign io_mops_ysyx_debug = 32'h6b == io_inst; // @[Decode.scala 387:35]
  assign io_mops_ysyx_print = 32'h7b == io_inst; // @[Decode.scala 388:35]
  assign io_mops_inst = io_inst; // @[Decode.scala 389:24]
endmodule
module Dec16(
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_bht_predict_taken,
  input  [31:0] io_target_pc,
  output        io_mops_illegal,
  output [3:0]  io_mops_next_pc,
  output [1:0]  io_mops_alu_mdu_lsu,
  output [3:0]  io_mops_branch_type,
  output [1:0]  io_mops_src_b,
  output        io_mops_write_dest,
  output [4:0]  io_mops_alu_op,
  output        io_mops_alu_expand,
  output [2:0]  io_mops_mem_width,
  output [1:0]  io_mops_write_src,
  output [4:0]  io_mops_rs1,
  output [4:0]  io_mops_rs2,
  output [4:0]  io_mops_rd,
  output [19:0] io_mops_imm,
  output [31:0] io_mops_pc,
  output        io_mops_predict_taken,
  output [31:0] io_mops_target_pc,
  output [31:0] io_mops_inst
);
  wire [31:0] _control_signal_T = io_inst & 32'he003; // @[Lookup.scala 31:38]
  wire  _control_signal_T_1 = 32'h0 == _control_signal_T; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_2 = io_inst & 32'hef83; // @[Lookup.scala 31:38]
  wire  _control_signal_T_3 = 32'h1 == _control_signal_T_2; // @[Lookup.scala 31:38]
  wire  _control_signal_T_5 = 32'h1 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_7 = 32'h2001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_9 = 32'h4001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_11 = 32'h6101 == _control_signal_T_2; // @[Lookup.scala 31:38]
  wire  _control_signal_T_13 = 32'h6001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_14 = io_inst & 32'hec03; // @[Lookup.scala 31:38]
  wire  _control_signal_T_15 = 32'h8001 == _control_signal_T_14; // @[Lookup.scala 31:38]
  wire  _control_signal_T_17 = 32'h8401 == _control_signal_T_14; // @[Lookup.scala 31:38]
  wire  _control_signal_T_19 = 32'h8801 == _control_signal_T_14; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_20 = io_inst & 32'hfc63; // @[Lookup.scala 31:38]
  wire  _control_signal_T_21 = 32'h8c01 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_23 = 32'h8c21 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_25 = 32'h8c41 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_27 = 32'h8c61 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_29 = 32'h9c01 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_31 = 32'h9c21 == _control_signal_T_20; // @[Lookup.scala 31:38]
  wire  _control_signal_T_33 = 32'h2 == _control_signal_T; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_34 = io_inst & 32'hf003; // @[Lookup.scala 31:38]
  wire  _control_signal_T_35 = 32'h8002 == _control_signal_T_34; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_36 = io_inst & 32'hffff; // @[Lookup.scala 31:38]
  wire  _control_signal_T_37 = 32'h9002 == _control_signal_T_36; // @[Lookup.scala 31:38]
  wire  _control_signal_T_39 = 32'h9002 == _control_signal_T_34; // @[Lookup.scala 31:38]
  wire  _control_signal_T_41 = 32'h4000 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_43 = 32'h6000 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_45 = 32'hc000 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_47 = 32'he000 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_49 = 32'h4002 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_51 = 32'h6002 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_53 = 32'hc002 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_55 = 32'he002 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_57 = 32'ha001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_59 = 32'hc001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire  _control_signal_T_61 = 32'he001 == _control_signal_T; // @[Lookup.scala 31:38]
  wire [31:0] _control_signal_T_62 = io_inst & 32'hf07f; // @[Lookup.scala 31:38]
  wire  _control_signal_T_63 = 32'h8002 == _control_signal_T_62; // @[Lookup.scala 31:38]
  wire  _control_signal_T_65 = 32'h9002 == _control_signal_T_62; // @[Lookup.scala 31:38]
  wire  _control_signal_T_66 = _control_signal_T_65 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  wire  _control_signal_T_67 = _control_signal_T_63 ? 1'h0 : _control_signal_T_66; // @[Lookup.scala 33:37]
  wire  _control_signal_T_68 = _control_signal_T_61 ? 1'h0 : _control_signal_T_67; // @[Lookup.scala 33:37]
  wire  _control_signal_T_69 = _control_signal_T_59 ? 1'h0 : _control_signal_T_68; // @[Lookup.scala 33:37]
  wire  _control_signal_T_70 = _control_signal_T_57 ? 1'h0 : _control_signal_T_69; // @[Lookup.scala 33:37]
  wire  _control_signal_T_71 = _control_signal_T_55 ? 1'h0 : _control_signal_T_70; // @[Lookup.scala 33:37]
  wire  _control_signal_T_72 = _control_signal_T_53 ? 1'h0 : _control_signal_T_71; // @[Lookup.scala 33:37]
  wire  _control_signal_T_73 = _control_signal_T_51 ? 1'h0 : _control_signal_T_72; // @[Lookup.scala 33:37]
  wire  _control_signal_T_74 = _control_signal_T_49 ? 1'h0 : _control_signal_T_73; // @[Lookup.scala 33:37]
  wire  _control_signal_T_75 = _control_signal_T_47 ? 1'h0 : _control_signal_T_74; // @[Lookup.scala 33:37]
  wire  _control_signal_T_76 = _control_signal_T_45 ? 1'h0 : _control_signal_T_75; // @[Lookup.scala 33:37]
  wire  _control_signal_T_77 = _control_signal_T_43 ? 1'h0 : _control_signal_T_76; // @[Lookup.scala 33:37]
  wire  _control_signal_T_78 = _control_signal_T_41 ? 1'h0 : _control_signal_T_77; // @[Lookup.scala 33:37]
  wire  _control_signal_T_79 = _control_signal_T_39 ? 1'h0 : _control_signal_T_78; // @[Lookup.scala 33:37]
  wire  _control_signal_T_80 = _control_signal_T_37 ? 1'h0 : _control_signal_T_79; // @[Lookup.scala 33:37]
  wire  _control_signal_T_81 = _control_signal_T_35 ? 1'h0 : _control_signal_T_80; // @[Lookup.scala 33:37]
  wire  _control_signal_T_82 = _control_signal_T_33 ? 1'h0 : _control_signal_T_81; // @[Lookup.scala 33:37]
  wire  _control_signal_T_83 = _control_signal_T_31 ? 1'h0 : _control_signal_T_82; // @[Lookup.scala 33:37]
  wire  _control_signal_T_84 = _control_signal_T_29 ? 1'h0 : _control_signal_T_83; // @[Lookup.scala 33:37]
  wire  _control_signal_T_85 = _control_signal_T_27 ? 1'h0 : _control_signal_T_84; // @[Lookup.scala 33:37]
  wire  _control_signal_T_86 = _control_signal_T_25 ? 1'h0 : _control_signal_T_85; // @[Lookup.scala 33:37]
  wire  _control_signal_T_87 = _control_signal_T_23 ? 1'h0 : _control_signal_T_86; // @[Lookup.scala 33:37]
  wire  _control_signal_T_88 = _control_signal_T_21 ? 1'h0 : _control_signal_T_87; // @[Lookup.scala 33:37]
  wire  _control_signal_T_89 = _control_signal_T_19 ? 1'h0 : _control_signal_T_88; // @[Lookup.scala 33:37]
  wire  _control_signal_T_90 = _control_signal_T_17 ? 1'h0 : _control_signal_T_89; // @[Lookup.scala 33:37]
  wire  _control_signal_T_91 = _control_signal_T_15 ? 1'h0 : _control_signal_T_90; // @[Lookup.scala 33:37]
  wire  _control_signal_T_92 = _control_signal_T_13 ? 1'h0 : _control_signal_T_91; // @[Lookup.scala 33:37]
  wire  _control_signal_T_93 = _control_signal_T_11 ? 1'h0 : _control_signal_T_92; // @[Lookup.scala 33:37]
  wire  _control_signal_T_94 = _control_signal_T_9 ? 1'h0 : _control_signal_T_93; // @[Lookup.scala 33:37]
  wire  _control_signal_T_95 = _control_signal_T_7 ? 1'h0 : _control_signal_T_94; // @[Lookup.scala 33:37]
  wire  _control_signal_T_96 = _control_signal_T_5 ? 1'h0 : _control_signal_T_95; // @[Lookup.scala 33:37]
  wire  _control_signal_T_97 = _control_signal_T_3 ? 1'h0 : _control_signal_T_96; // @[Lookup.scala 33:37]
  wire  control_signal_0 = _control_signal_T_1 ? 1'h0 : _control_signal_T_97; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_103 = _control_signal_T_55 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_104 = _control_signal_T_53 ? 2'h2 : _control_signal_T_103; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_105 = _control_signal_T_51 ? 2'h2 : _control_signal_T_104; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_106 = _control_signal_T_49 ? 2'h2 : _control_signal_T_105; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_107 = _control_signal_T_47 ? 2'h2 : _control_signal_T_106; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_108 = _control_signal_T_45 ? 2'h2 : _control_signal_T_107; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_109 = _control_signal_T_43 ? 2'h2 : _control_signal_T_108; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_110 = _control_signal_T_41 ? 2'h2 : _control_signal_T_109; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_111 = _control_signal_T_39 ? 2'h3 : _control_signal_T_110; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_112 = _control_signal_T_37 ? 2'h0 : _control_signal_T_111; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_113 = _control_signal_T_35 ? 2'h3 : _control_signal_T_112; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_114 = _control_signal_T_33 ? 2'h3 : _control_signal_T_113; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_115 = _control_signal_T_31 ? 2'h3 : _control_signal_T_114; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_116 = _control_signal_T_29 ? 2'h3 : _control_signal_T_115; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_117 = _control_signal_T_27 ? 2'h3 : _control_signal_T_116; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_118 = _control_signal_T_25 ? 2'h3 : _control_signal_T_117; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_119 = _control_signal_T_23 ? 2'h3 : _control_signal_T_118; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_120 = _control_signal_T_21 ? 2'h3 : _control_signal_T_119; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_121 = _control_signal_T_19 ? 2'h3 : _control_signal_T_120; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_122 = _control_signal_T_17 ? 2'h3 : _control_signal_T_121; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_123 = _control_signal_T_15 ? 2'h3 : _control_signal_T_122; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_124 = _control_signal_T_13 ? 2'h3 : _control_signal_T_123; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_125 = _control_signal_T_11 ? 2'h3 : _control_signal_T_124; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_126 = _control_signal_T_9 ? 2'h3 : _control_signal_T_125; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_127 = _control_signal_T_7 ? 2'h3 : _control_signal_T_126; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_128 = _control_signal_T_5 ? 2'h3 : _control_signal_T_127; // @[Lookup.scala 33:37]
  wire [1:0] _control_signal_T_129 = _control_signal_T_3 ? 2'h3 : _control_signal_T_128; // @[Lookup.scala 33:37]
  wire [1:0] control_signal_1 = _control_signal_T_1 ? 2'h3 : _control_signal_T_129; // @[Lookup.scala 33:37]
  wire [4:0] CREG1 = io_inst[11:7]; // @[Decode.scala 453:24]
  wire [4:0] CREG2 = io_inst[6:2]; // @[Decode.scala 454:24]
  wire [2:0] CREG1P_lo = io_inst[4:2]; // @[Decode.scala 455:32]
  wire [4:0] CREG1P = {2'h1,CREG1P_lo}; // @[Cat.scala 30:58]
  wire [2:0] CREG2P_lo = io_inst[9:7]; // @[Decode.scala 456:32]
  wire [4:0] CREG2P = {2'h1,CREG2P_lo}; // @[Cat.scala 30:58]
  wire [14:0] IIMM_hi = io_inst[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [19:0] IIMM = {IIMM_hi,CREG2}; // @[Cat.scala 30:58]
  wire [2:0] LUIIMM_hi_hi = io_inst[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [19:0] LUIIMM = {LUIIMM_hi_hi,CREG2,12'h0}; // @[Cat.scala 30:58]
  wire [10:0] ADDI16SPIMM_hi_hi = io_inst[12] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [19:0] ADDI16SPIMM = {ADDI16SPIMM_hi_hi,CREG2,4'h0}; // @[Cat.scala 30:58]
  wire [3:0] ADDI4SPNIMM_hi_hi_lo = io_inst[10:7]; // @[Decode.scala 463:56]
  wire [1:0] ADDI4SPNIMM_hi_lo = io_inst[12:11]; // @[Decode.scala 463:72]
  wire  ADDI4SPNIMM_lo_hi_hi = io_inst[5]; // @[Decode.scala 463:89]
  wire  ADDI4SPNIMM_lo_hi_lo = io_inst[6]; // @[Decode.scala 463:101]
  wire [19:0] ADDI4SPNIMM = {10'h0,ADDI4SPNIMM_hi_hi_lo,ADDI4SPNIMM_hi_lo,ADDI4SPNIMM_lo_hi_hi,ADDI4SPNIMM_lo_hi_lo,2'h0
    }; // @[Cat.scala 30:58]
  wire [19:0] SHAMT = {14'h0,io_inst[12],CREG2}; // @[Cat.scala 30:58]
  wire [4:0] _alu_signal_T_39 = _control_signal_T_29 ? CREG2P : CREG1; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_40 = _control_signal_T_31 ? CREG2P : _alu_signal_T_39; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_41 = _control_signal_T_21 ? CREG2P : _alu_signal_T_40; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_42 = _control_signal_T_23 ? CREG2P : _alu_signal_T_41; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_43 = _control_signal_T_25 ? CREG2P : _alu_signal_T_42; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_44 = _control_signal_T_27 ? CREG2P : _alu_signal_T_43; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_45 = _control_signal_T_39 ? CREG1 : _alu_signal_T_44; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_46 = _control_signal_T_35 ? CREG1 : _alu_signal_T_45; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_47 = _control_signal_T_19 ? CREG2P : _alu_signal_T_46; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_48 = _control_signal_T_17 ? CREG2P : _alu_signal_T_47; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_49 = _control_signal_T_15 ? CREG2P : _alu_signal_T_48; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_50 = _control_signal_T_33 ? CREG1 : _alu_signal_T_49; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_51 = _control_signal_T_1 ? CREG1P : _alu_signal_T_50; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_52 = _control_signal_T_11 ? CREG1 : _alu_signal_T_51; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_53 = _control_signal_T_7 ? CREG1 : _alu_signal_T_52; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_54 = _control_signal_T_5 ? CREG1 : _alu_signal_T_53; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_55 = _control_signal_T_13 ? CREG1 : _alu_signal_T_54; // @[Lookup.scala 33:37]
  wire [4:0] alu_signal_0 = _control_signal_T_9 ? CREG1 : _alu_signal_T_55; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_64 = _control_signal_T_35 ? CREG2 : _alu_signal_T_45; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_65 = _control_signal_T_19 ? CREG2P : _alu_signal_T_64; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_66 = _control_signal_T_17 ? CREG2P : _alu_signal_T_65; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_67 = _control_signal_T_15 ? CREG2P : _alu_signal_T_66; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_68 = _control_signal_T_33 ? CREG1 : _alu_signal_T_67; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_69 = _control_signal_T_1 ? 5'h2 : _alu_signal_T_68; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_70 = _control_signal_T_11 ? CREG1 : _alu_signal_T_69; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_71 = _control_signal_T_7 ? CREG1 : _alu_signal_T_70; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_72 = _control_signal_T_5 ? CREG1 : _alu_signal_T_71; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_73 = _control_signal_T_13 ? 5'h0 : _alu_signal_T_72; // @[Lookup.scala 33:37]
  wire [4:0] alu_signal_1 = _control_signal_T_9 ? 5'h0 : _alu_signal_T_73; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_74 = _control_signal_T_3 ? 5'h0 : CREG2; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_75 = _control_signal_T_29 ? CREG1P : _alu_signal_T_74; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_76 = _control_signal_T_31 ? CREG1P : _alu_signal_T_75; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_77 = _control_signal_T_21 ? CREG1P : _alu_signal_T_76; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_78 = _control_signal_T_23 ? CREG1P : _alu_signal_T_77; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_79 = _control_signal_T_25 ? CREG1P : _alu_signal_T_78; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_80 = _control_signal_T_27 ? CREG1P : _alu_signal_T_79; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_81 = _control_signal_T_39 ? CREG2 : _alu_signal_T_80; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_82 = _control_signal_T_35 ? 5'h0 : _alu_signal_T_81; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_83 = _control_signal_T_19 ? 5'h0 : _alu_signal_T_82; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_84 = _control_signal_T_17 ? 5'h0 : _alu_signal_T_83; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_85 = _control_signal_T_15 ? 5'h0 : _alu_signal_T_84; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_86 = _control_signal_T_33 ? 5'h0 : _alu_signal_T_85; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_87 = _control_signal_T_1 ? 5'h0 : _alu_signal_T_86; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_88 = _control_signal_T_11 ? 5'h0 : _alu_signal_T_87; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_89 = _control_signal_T_7 ? 5'h0 : _alu_signal_T_88; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_90 = _control_signal_T_5 ? 5'h0 : _alu_signal_T_89; // @[Lookup.scala 33:37]
  wire [4:0] _alu_signal_T_91 = _control_signal_T_13 ? 5'h0 : _alu_signal_T_90; // @[Lookup.scala 33:37]
  wire [4:0] alu_signal_2 = _control_signal_T_9 ? 5'h0 : _alu_signal_T_91; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_101 = _control_signal_T_19 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_102 = _control_signal_T_17 ? 2'h1 : _alu_signal_T_101; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_103 = _control_signal_T_15 ? 2'h1 : _alu_signal_T_102; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_104 = _control_signal_T_33 ? 2'h1 : _alu_signal_T_103; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_105 = _control_signal_T_1 ? 2'h1 : _alu_signal_T_104; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_106 = _control_signal_T_11 ? 2'h1 : _alu_signal_T_105; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_107 = _control_signal_T_7 ? 2'h1 : _alu_signal_T_106; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_108 = _control_signal_T_5 ? 2'h1 : _alu_signal_T_107; // @[Lookup.scala 33:37]
  wire [1:0] _alu_signal_T_109 = _control_signal_T_13 ? 2'h1 : _alu_signal_T_108; // @[Lookup.scala 33:37]
  wire [1:0] alu_signal_3 = _control_signal_T_9 ? 2'h1 : _alu_signal_T_109; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_112 = _control_signal_T_31 ? 1'h0 : _control_signal_T_29; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_113 = _control_signal_T_21 | _alu_signal_T_112; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_114 = _control_signal_T_23 ? 3'h4 : {{2'd0}, _alu_signal_T_113}; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_115 = _control_signal_T_25 ? 3'h6 : _alu_signal_T_114; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_116 = _control_signal_T_27 ? 3'h5 : _alu_signal_T_115; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_117 = _control_signal_T_39 ? 3'h0 : _alu_signal_T_116; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_118 = _control_signal_T_35 ? 3'h0 : _alu_signal_T_117; // @[Lookup.scala 33:37]
  wire [2:0] _alu_signal_T_119 = _control_signal_T_19 ? 3'h5 : _alu_signal_T_118; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_120 = _control_signal_T_17 ? 4'h9 : {{1'd0}, _alu_signal_T_119}; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_121 = _control_signal_T_15 ? 4'h8 : _alu_signal_T_120; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_122 = _control_signal_T_33 ? 4'h7 : _alu_signal_T_121; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_123 = _control_signal_T_1 ? 4'h0 : _alu_signal_T_122; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_124 = _control_signal_T_11 ? 4'h0 : _alu_signal_T_123; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_125 = _control_signal_T_7 ? 4'h0 : _alu_signal_T_124; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_126 = _control_signal_T_5 ? 4'h0 : _alu_signal_T_125; // @[Lookup.scala 33:37]
  wire [3:0] _alu_signal_T_127 = _control_signal_T_13 ? 4'ha : _alu_signal_T_126; // @[Lookup.scala 33:37]
  wire [3:0] alu_signal_4 = _control_signal_T_9 ? 4'h0 : _alu_signal_T_127; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_137 = _control_signal_T_19 ? IIMM : 20'h0; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_138 = _control_signal_T_17 ? SHAMT : _alu_signal_T_137; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_139 = _control_signal_T_15 ? SHAMT : _alu_signal_T_138; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_140 = _control_signal_T_33 ? SHAMT : _alu_signal_T_139; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_141 = _control_signal_T_1 ? ADDI4SPNIMM : _alu_signal_T_140; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_142 = _control_signal_T_11 ? ADDI16SPIMM : _alu_signal_T_141; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_143 = _control_signal_T_7 ? IIMM : _alu_signal_T_142; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_144 = _control_signal_T_5 ? IIMM : _alu_signal_T_143; // @[Lookup.scala 33:37]
  wire [19:0] _alu_signal_T_145 = _control_signal_T_13 ? LUIIMM : _alu_signal_T_144; // @[Lookup.scala 33:37]
  wire [19:0] alu_signal_5 = _control_signal_T_9 ? IIMM : _alu_signal_T_145; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_149 = _control_signal_T_21 ? 1'h0 : _control_signal_T_31 | _control_signal_T_29; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_150 = _control_signal_T_23 ? 1'h0 : _alu_signal_T_149; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_151 = _control_signal_T_25 ? 1'h0 : _alu_signal_T_150; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_152 = _control_signal_T_27 ? 1'h0 : _alu_signal_T_151; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_153 = _control_signal_T_39 ? 1'h0 : _alu_signal_T_152; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_154 = _control_signal_T_35 ? 1'h0 : _alu_signal_T_153; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_155 = _control_signal_T_19 ? 1'h0 : _alu_signal_T_154; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_156 = _control_signal_T_17 ? 1'h0 : _alu_signal_T_155; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_157 = _control_signal_T_15 ? 1'h0 : _alu_signal_T_156; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_158 = _control_signal_T_33 ? 1'h0 : _alu_signal_T_157; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_159 = _control_signal_T_1 ? 1'h0 : _alu_signal_T_158; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_160 = _control_signal_T_11 ? 1'h0 : _alu_signal_T_159; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_162 = _control_signal_T_5 ? 1'h0 : _control_signal_T_7 | _alu_signal_T_160; // @[Lookup.scala 33:37]
  wire  _alu_signal_T_163 = _control_signal_T_13 ? 1'h0 : _alu_signal_T_162; // @[Lookup.scala 33:37]
  wire  alu_signal_6 = _control_signal_T_9 ? 1'h0 : _alu_signal_T_163; // @[Lookup.scala 33:37]
  wire [1:0] LWSPIMM_hi_lo = io_inst[3:2]; // @[Decode.scala 492:39]
  wire [2:0] LWSPIMM_lo_hi = io_inst[6:4]; // @[Decode.scala 492:54]
  wire [62:0] LWSPIMM = {56'h0,LWSPIMM_hi_lo,LWSPIMM_lo_hi,2'h0}; // @[Cat.scala 30:58]
  wire [1:0] LDSPIMM_lo_hi = io_inst[6:5]; // @[Decode.scala 493:54]
  wire [62:0] LDSPIMM = {55'h0,CREG1P_lo,LDSPIMM_lo_hi,3'h0}; // @[Cat.scala 30:58]
  wire [1:0] SWSPIMM_hi_lo = io_inst[8:7]; // @[Decode.scala 494:39]
  wire [3:0] SWSPIMM_lo_hi = io_inst[12:9]; // @[Decode.scala 494:54]
  wire [63:0] SWSPIMM = {56'h0,SWSPIMM_hi_lo,SWSPIMM_lo_hi,2'h0}; // @[Cat.scala 30:58]
  wire [2:0] SDSPIMM_lo_hi = io_inst[12:10]; // @[Decode.scala 495:54]
  wire [63:0] SDSPIMM = {55'h0,CREG2P_lo,SDSPIMM_lo_hi,3'h0}; // @[Cat.scala 30:58]
  wire [63:0] WIMM = {57'h0,ADDI4SPNIMM_lo_hi_hi,SDSPIMM_lo_hi,ADDI4SPNIMM_lo_hi_lo,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] DIMM = {56'h0,LDSPIMM_lo_hi,SDSPIMM_lo_hi,3'h0}; // @[Cat.scala 30:58]
  wire [4:0] _lsu_signal_T_16 = _control_signal_T_45 ? 5'h0 : CREG1P; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_17 = _control_signal_T_45 ? 5'h0 : _lsu_signal_T_16; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_18 = _control_signal_T_43 ? CREG1P : _lsu_signal_T_17; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_19 = _control_signal_T_41 ? CREG1P : _lsu_signal_T_18; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_20 = _control_signal_T_55 ? 5'h0 : _lsu_signal_T_19; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_21 = _control_signal_T_53 ? 5'h0 : _lsu_signal_T_20; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_22 = _control_signal_T_51 ? CREG1 : _lsu_signal_T_21; // @[Lookup.scala 33:37]
  wire [4:0] lsu_signal_0 = _control_signal_T_49 ? CREG1 : _lsu_signal_T_22; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_27 = _control_signal_T_55 ? 5'h2 : CREG2P; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_28 = _control_signal_T_53 ? 5'h2 : _lsu_signal_T_27; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_29 = _control_signal_T_51 ? 5'h2 : _lsu_signal_T_28; // @[Lookup.scala 33:37]
  wire [4:0] lsu_signal_1 = _control_signal_T_49 ? 5'h2 : _lsu_signal_T_29; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_30 = _control_signal_T_45 ? CREG1P : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_31 = _control_signal_T_45 ? CREG1P : _lsu_signal_T_30; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_32 = _control_signal_T_43 ? 5'h0 : _lsu_signal_T_31; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_33 = _control_signal_T_41 ? 5'h0 : _lsu_signal_T_32; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_34 = _control_signal_T_55 ? CREG2 : _lsu_signal_T_33; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_35 = _control_signal_T_53 ? CREG2 : _lsu_signal_T_34; // @[Lookup.scala 33:37]
  wire [4:0] _lsu_signal_T_36 = _control_signal_T_51 ? 5'h0 : _lsu_signal_T_35; // @[Lookup.scala 33:37]
  wire [4:0] lsu_signal_2 = _control_signal_T_49 ? 5'h0 : _lsu_signal_T_36; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_37 = _control_signal_T_45 ? DIMM : WIMM; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_38 = _control_signal_T_45 ? WIMM : _lsu_signal_T_37; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_39 = _control_signal_T_43 ? DIMM : _lsu_signal_T_38; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_40 = _control_signal_T_41 ? WIMM : _lsu_signal_T_39; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_41 = _control_signal_T_55 ? SDSPIMM : _lsu_signal_T_40; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_42 = _control_signal_T_53 ? SWSPIMM : _lsu_signal_T_41; // @[Lookup.scala 33:37]
  wire [63:0] _lsu_signal_T_43 = _control_signal_T_51 ? {{1'd0}, LDSPIMM} : _lsu_signal_T_42; // @[Lookup.scala 33:37]
  wire [63:0] lsu_signal_3 = _control_signal_T_49 ? {{1'd0}, LWSPIMM} : _lsu_signal_T_43; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_44 = _control_signal_T_45 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_45 = _control_signal_T_45 ? 1'h0 : _lsu_signal_T_44; // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_48 = _control_signal_T_55 ? 1'h0 : _control_signal_T_41 | (_control_signal_T_43 | _lsu_signal_T_45
    ); // @[Lookup.scala 33:37]
  wire  _lsu_signal_T_49 = _control_signal_T_53 ? 1'h0 : _lsu_signal_T_48; // @[Lookup.scala 33:37]
  wire  lsu_signal_4 = _control_signal_T_49 | (_control_signal_T_51 | _lsu_signal_T_49); // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_51 = _control_signal_T_45 ? 3'h5 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_52 = _control_signal_T_45 ? 3'h4 : _lsu_signal_T_51; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_53 = _control_signal_T_43 ? 3'h5 : _lsu_signal_T_52; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_54 = _control_signal_T_41 ? 3'h4 : _lsu_signal_T_53; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_55 = _control_signal_T_55 ? 3'h5 : _lsu_signal_T_54; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_56 = _control_signal_T_53 ? 3'h4 : _lsu_signal_T_55; // @[Lookup.scala 33:37]
  wire [2:0] _lsu_signal_T_57 = _control_signal_T_51 ? 3'h5 : _lsu_signal_T_56; // @[Lookup.scala 33:37]
  wire [2:0] lsu_signal_5 = _control_signal_T_49 ? 3'h4 : _lsu_signal_T_57; // @[Lookup.scala 33:37]
  wire [55:0] BIMM_hi_hi_hi = io_inst[12] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire  BIMM_hi_lo = io_inst[2]; // @[Decode.scala 512:64]
  wire [1:0] BIMM_lo_hi_hi = io_inst[11:10]; // @[Decode.scala 512:76]
  wire [1:0] BIMM_lo_hi_lo = io_inst[4:3]; // @[Decode.scala 512:93]
  wire [63:0] BIMM = {BIMM_hi_hi_hi,LDSPIMM_lo_hi,BIMM_hi_lo,BIMM_lo_hi_hi,BIMM_lo_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [52:0] JIMM_hi_hi_hi_hi = io_inst[12] ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  wire  JIMM_hi_hi_hi_lo = io_inst[8]; // @[Decode.scala 513:49]
  wire [1:0] JIMM_hi_hi_lo = io_inst[10:9]; // @[Decode.scala 513:61]
  wire  JIMM_hi_lo_lo = io_inst[7]; // @[Decode.scala 513:89]
  wire  JIMM_lo_hi_lo = io_inst[11]; // @[Decode.scala 513:113]
  wire [2:0] JIMM_lo_lo_hi = io_inst[5:3]; // @[Decode.scala 513:126]
  wire [63:0] JIMM = {JIMM_hi_hi_hi_hi,JIMM_hi_hi_hi_lo,JIMM_hi_hi_lo,ADDI4SPNIMM_lo_hi_lo,JIMM_hi_lo_lo,BIMM_hi_lo,
    JIMM_lo_hi_lo,JIMM_lo_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [3:0] _bju_signal_T_10 = _control_signal_T_61 ? 4'h2 : 4'h1; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_11 = _control_signal_T_59 ? 4'h2 : _bju_signal_T_10; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_12 = _control_signal_T_65 ? 4'h4 : _bju_signal_T_11; // @[Lookup.scala 33:37]
  wire [3:0] _bju_signal_T_13 = _control_signal_T_63 ? 4'h4 : _bju_signal_T_12; // @[Lookup.scala 33:37]
  wire [3:0] bju_signal_0 = _control_signal_T_57 ? 4'h3 : _bju_signal_T_13; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_14 = _control_signal_T_61 ? CREG2P : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_15 = _control_signal_T_59 ? CREG2P : _bju_signal_T_14; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_16 = _control_signal_T_65 ? 5'h1 : _bju_signal_T_15; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_17 = _control_signal_T_63 ? 5'h0 : _bju_signal_T_16; // @[Lookup.scala 33:37]
  wire [4:0] bju_signal_1 = _control_signal_T_57 ? 5'h0 : _bju_signal_T_17; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_20 = _control_signal_T_65 ? CREG1 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _bju_signal_T_21 = _control_signal_T_63 ? CREG1 : _bju_signal_T_20; // @[Lookup.scala 33:37]
  wire [4:0] bju_signal_2 = _control_signal_T_57 ? 5'h0 : _bju_signal_T_21; // @[Lookup.scala 33:37]
  wire  bju_signal_4 = _control_signal_T_57 | (_control_signal_T_63 | _control_signal_T_65); // @[Lookup.scala 33:37]
  wire  _bju_signal_T_32 = _control_signal_T_65 ? 1'h0 : _control_signal_T_59 | _control_signal_T_61; // @[Lookup.scala 33:37]
  wire  _bju_signal_T_33 = _control_signal_T_63 ? 1'h0 : _bju_signal_T_32; // @[Lookup.scala 33:37]
  wire  bju_signal_5 = _control_signal_T_57 ? 1'h0 : _bju_signal_T_33; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_34 = _control_signal_T_61 ? BIMM : 64'h0; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_35 = _control_signal_T_59 ? BIMM : _bju_signal_T_34; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_36 = _control_signal_T_65 ? 64'h0 : _bju_signal_T_35; // @[Lookup.scala 33:37]
  wire [63:0] _bju_signal_T_37 = _control_signal_T_63 ? 64'h0 : _bju_signal_T_36; // @[Lookup.scala 33:37]
  wire [63:0] bju_signal_6 = _control_signal_T_57 ? JIMM : _bju_signal_T_37; // @[Lookup.scala 33:37]
  wire [3:0] branch_signal_0 = _control_signal_T_59 ? 4'h1 : _bju_signal_T_10; // @[Lookup.scala 33:37]
  wire  _io_mops_branch_type_T = control_signal_1 == 2'h0; // @[Decode.scala 541:50]
  wire  _io_mops_src_b_T = control_signal_1 == 2'h3; // @[Decode.scala 545:50]
  wire  _io_mops_write_dest_T_1 = 2'h2 == control_signal_1 ? lsu_signal_4 : 1'h1; // @[Mux.scala 80:57]
  wire [3:0] _io_mops_alu_op_T_1 = 2'h3 == control_signal_1 ? alu_signal_4 : 4'h0; // @[Mux.scala 80:57]
  wire [3:0] _io_mops_alu_op_T_3 = 2'h0 == control_signal_1 ? {{3'd0}, bju_signal_5} : _io_mops_alu_op_T_1; // @[Mux.scala 80:57]
  wire [1:0] _io_mops_write_src_T_3 = bju_signal_0 == 4'h3 | bju_signal_0 == 4'h4 ? 2'h3 : 2'h0; // @[Decode.scala 563:21]
  wire [1:0] _io_mops_write_src_T_5 = 2'h2 == control_signal_1 ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs1_T_1 = 2'h2 == control_signal_1 ? lsu_signal_1 : alu_signal_1; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rs2_T_1 = 2'h2 == control_signal_1 ? lsu_signal_2 : alu_signal_2; // @[Mux.scala 80:57]
  wire [4:0] _io_mops_rd_T_1 = 2'h2 == control_signal_1 ? lsu_signal_0 : alu_signal_0; // @[Mux.scala 80:57]
  wire [63:0] _io_mops_imm_T_1 = 2'h2 == control_signal_1 ? lsu_signal_3 : {{44'd0}, alu_signal_5}; // @[Mux.scala 80:57]
  wire [63:0] _io_mops_imm_T_3 = 2'h0 == control_signal_1 ? bju_signal_6 : _io_mops_imm_T_1; // @[Mux.scala 80:57]
  wire [47:0] _io_mops_inst_T = {16'h0,io_inst}; // @[Cat.scala 30:58]
  assign io_mops_illegal = control_signal_0 | |io_pc[1:0]; // @[Decode.scala 540:53]
  assign io_mops_next_pc = _io_mops_branch_type_T ? bju_signal_0 : 4'h1; // @[Decode.scala 543:31]
  assign io_mops_alu_mdu_lsu = _control_signal_T_1 ? 2'h3 : _control_signal_T_129; // @[Lookup.scala 33:37]
  assign io_mops_branch_type = control_signal_1 == 2'h0 & bju_signal_0 == 4'h2 ? branch_signal_0 : 4'h0; // @[Decode.scala 541:31]
  assign io_mops_src_b = control_signal_1 == 2'h3 ? alu_signal_3 : 2'h1; // @[Decode.scala 545:31]
  assign io_mops_write_dest = 2'h0 == control_signal_1 ? bju_signal_4 : _io_mops_write_dest_T_1; // @[Mux.scala 80:57]
  assign io_mops_alu_op = {{1'd0}, _io_mops_alu_op_T_3}; // @[Mux.scala 80:57]
  assign io_mops_alu_expand = _io_mops_src_b_T & alu_signal_6; // @[Decode.scala 558:31]
  assign io_mops_mem_width = control_signal_1 == 2'h2 ? lsu_signal_5 : 3'h0; // @[Decode.scala 559:31]
  assign io_mops_write_src = 2'h0 == control_signal_1 ? _io_mops_write_src_T_3 : _io_mops_write_src_T_5; // @[Mux.scala 80:57]
  assign io_mops_rs1 = 2'h0 == control_signal_1 ? bju_signal_1 : _io_mops_rs1_T_1; // @[Mux.scala 80:57]
  assign io_mops_rs2 = 2'h0 == control_signal_1 ? bju_signal_2 : _io_mops_rs2_T_1; // @[Mux.scala 80:57]
  assign io_mops_rd = 2'h0 == control_signal_1 ? 5'h0 : _io_mops_rd_T_1; // @[Mux.scala 80:57]
  assign io_mops_imm = _io_mops_imm_T_3[19:0]; // @[Decode.scala 584:25]
  assign io_mops_pc = io_pc; // @[Decode.scala 590:25]
  assign io_mops_predict_taken = io_bht_predict_taken; // @[Decode.scala 591:25]
  assign io_mops_target_pc = io_target_pc; // @[Decode.scala 592:25]
  assign io_mops_inst = _io_mops_inst_T[31:0]; // @[Decode.scala 596:24]
endmodule
module Dec(
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_bht_predict_taken,
  input  [31:0] io_target_pc,
  output        io_mops_illegal,
  output [3:0]  io_mops_next_pc,
  output [1:0]  io_mops_alu_mdu_lsu,
  output [3:0]  io_mops_branch_type,
  output [1:0]  io_mops_src_a,
  output [1:0]  io_mops_src_b,
  output        io_mops_write_dest,
  output [4:0]  io_mops_alu_op,
  output        io_mops_alu_expand,
  output [2:0]  io_mops_mem_width,
  output [1:0]  io_mops_write_src,
  output [4:0]  io_mops_rs1,
  output [4:0]  io_mops_rs2,
  output [4:0]  io_mops_rd,
  output [19:0] io_mops_imm,
  output [31:0] io_mops_pc,
  output        io_mops_predict_taken,
  output [31:0] io_mops_target_pc,
  output        io_mops_ysyx_debug,
  output        io_mops_ysyx_print,
  output [31:0] io_mops_inst
);
  wire [31:0] decoder32_io_pc; // @[Decode.scala 46:25]
  wire [31:0] decoder32_io_inst; // @[Decode.scala 46:25]
  wire  decoder32_io_bht_predict_taken; // @[Decode.scala 46:25]
  wire [31:0] decoder32_io_target_pc; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_illegal; // @[Decode.scala 46:25]
  wire [3:0] decoder32_io_mops_next_pc; // @[Decode.scala 46:25]
  wire [1:0] decoder32_io_mops_alu_mdu_lsu; // @[Decode.scala 46:25]
  wire [3:0] decoder32_io_mops_branch_type; // @[Decode.scala 46:25]
  wire [1:0] decoder32_io_mops_src_a; // @[Decode.scala 46:25]
  wire [1:0] decoder32_io_mops_src_b; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_write_dest; // @[Decode.scala 46:25]
  wire [4:0] decoder32_io_mops_alu_op; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_alu_expand; // @[Decode.scala 46:25]
  wire [2:0] decoder32_io_mops_mem_width; // @[Decode.scala 46:25]
  wire [1:0] decoder32_io_mops_write_src; // @[Decode.scala 46:25]
  wire [4:0] decoder32_io_mops_rs1; // @[Decode.scala 46:25]
  wire [4:0] decoder32_io_mops_rs2; // @[Decode.scala 46:25]
  wire [4:0] decoder32_io_mops_rd; // @[Decode.scala 46:25]
  wire [19:0] decoder32_io_mops_imm; // @[Decode.scala 46:25]
  wire [31:0] decoder32_io_mops_pc; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_predict_taken; // @[Decode.scala 46:25]
  wire [31:0] decoder32_io_mops_target_pc; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_ysyx_debug; // @[Decode.scala 46:25]
  wire  decoder32_io_mops_ysyx_print; // @[Decode.scala 46:25]
  wire [31:0] decoder32_io_mops_inst; // @[Decode.scala 46:25]
  wire [31:0] decoder16_io_pc; // @[Decode.scala 47:25]
  wire [31:0] decoder16_io_inst; // @[Decode.scala 47:25]
  wire  decoder16_io_bht_predict_taken; // @[Decode.scala 47:25]
  wire [31:0] decoder16_io_target_pc; // @[Decode.scala 47:25]
  wire  decoder16_io_mops_illegal; // @[Decode.scala 47:25]
  wire [3:0] decoder16_io_mops_next_pc; // @[Decode.scala 47:25]
  wire [1:0] decoder16_io_mops_alu_mdu_lsu; // @[Decode.scala 47:25]
  wire [3:0] decoder16_io_mops_branch_type; // @[Decode.scala 47:25]
  wire [1:0] decoder16_io_mops_src_b; // @[Decode.scala 47:25]
  wire  decoder16_io_mops_write_dest; // @[Decode.scala 47:25]
  wire [4:0] decoder16_io_mops_alu_op; // @[Decode.scala 47:25]
  wire  decoder16_io_mops_alu_expand; // @[Decode.scala 47:25]
  wire [2:0] decoder16_io_mops_mem_width; // @[Decode.scala 47:25]
  wire [1:0] decoder16_io_mops_write_src; // @[Decode.scala 47:25]
  wire [4:0] decoder16_io_mops_rs1; // @[Decode.scala 47:25]
  wire [4:0] decoder16_io_mops_rs2; // @[Decode.scala 47:25]
  wire [4:0] decoder16_io_mops_rd; // @[Decode.scala 47:25]
  wire [19:0] decoder16_io_mops_imm; // @[Decode.scala 47:25]
  wire [31:0] decoder16_io_mops_pc; // @[Decode.scala 47:25]
  wire  decoder16_io_mops_predict_taken; // @[Decode.scala 47:25]
  wire [31:0] decoder16_io_mops_target_pc; // @[Decode.scala 47:25]
  wire [31:0] decoder16_io_mops_inst; // @[Decode.scala 47:25]
  Dec32 decoder32 ( // @[Decode.scala 46:25]
    .io_pc(decoder32_io_pc),
    .io_inst(decoder32_io_inst),
    .io_bht_predict_taken(decoder32_io_bht_predict_taken),
    .io_target_pc(decoder32_io_target_pc),
    .io_mops_illegal(decoder32_io_mops_illegal),
    .io_mops_next_pc(decoder32_io_mops_next_pc),
    .io_mops_alu_mdu_lsu(decoder32_io_mops_alu_mdu_lsu),
    .io_mops_branch_type(decoder32_io_mops_branch_type),
    .io_mops_src_a(decoder32_io_mops_src_a),
    .io_mops_src_b(decoder32_io_mops_src_b),
    .io_mops_write_dest(decoder32_io_mops_write_dest),
    .io_mops_alu_op(decoder32_io_mops_alu_op),
    .io_mops_alu_expand(decoder32_io_mops_alu_expand),
    .io_mops_mem_width(decoder32_io_mops_mem_width),
    .io_mops_write_src(decoder32_io_mops_write_src),
    .io_mops_rs1(decoder32_io_mops_rs1),
    .io_mops_rs2(decoder32_io_mops_rs2),
    .io_mops_rd(decoder32_io_mops_rd),
    .io_mops_imm(decoder32_io_mops_imm),
    .io_mops_pc(decoder32_io_mops_pc),
    .io_mops_predict_taken(decoder32_io_mops_predict_taken),
    .io_mops_target_pc(decoder32_io_mops_target_pc),
    .io_mops_ysyx_debug(decoder32_io_mops_ysyx_debug),
    .io_mops_ysyx_print(decoder32_io_mops_ysyx_print),
    .io_mops_inst(decoder32_io_mops_inst)
  );
  Dec16 decoder16 ( // @[Decode.scala 47:25]
    .io_pc(decoder16_io_pc),
    .io_inst(decoder16_io_inst),
    .io_bht_predict_taken(decoder16_io_bht_predict_taken),
    .io_target_pc(decoder16_io_target_pc),
    .io_mops_illegal(decoder16_io_mops_illegal),
    .io_mops_next_pc(decoder16_io_mops_next_pc),
    .io_mops_alu_mdu_lsu(decoder16_io_mops_alu_mdu_lsu),
    .io_mops_branch_type(decoder16_io_mops_branch_type),
    .io_mops_src_b(decoder16_io_mops_src_b),
    .io_mops_write_dest(decoder16_io_mops_write_dest),
    .io_mops_alu_op(decoder16_io_mops_alu_op),
    .io_mops_alu_expand(decoder16_io_mops_alu_expand),
    .io_mops_mem_width(decoder16_io_mops_mem_width),
    .io_mops_write_src(decoder16_io_mops_write_src),
    .io_mops_rs1(decoder16_io_mops_rs1),
    .io_mops_rs2(decoder16_io_mops_rs2),
    .io_mops_rd(decoder16_io_mops_rd),
    .io_mops_imm(decoder16_io_mops_imm),
    .io_mops_pc(decoder16_io_mops_pc),
    .io_mops_predict_taken(decoder16_io_mops_predict_taken),
    .io_mops_target_pc(decoder16_io_mops_target_pc),
    .io_mops_inst(decoder16_io_mops_inst)
  );
  assign io_mops_illegal = io_inst[1:0] == 2'h3 ? decoder32_io_mops_illegal : decoder16_io_mops_illegal; // @[Decode.scala 59:17]
  assign io_mops_next_pc = io_inst[1:0] == 2'h3 ? decoder32_io_mops_next_pc : decoder16_io_mops_next_pc; // @[Decode.scala 59:17]
  assign io_mops_alu_mdu_lsu = io_inst[1:0] == 2'h3 ? decoder32_io_mops_alu_mdu_lsu : decoder16_io_mops_alu_mdu_lsu; // @[Decode.scala 59:17]
  assign io_mops_branch_type = io_inst[1:0] == 2'h3 ? decoder32_io_mops_branch_type : decoder16_io_mops_branch_type; // @[Decode.scala 59:17]
  assign io_mops_src_a = io_inst[1:0] == 2'h3 ? decoder32_io_mops_src_a : 2'h0; // @[Decode.scala 59:17]
  assign io_mops_src_b = io_inst[1:0] == 2'h3 ? decoder32_io_mops_src_b : decoder16_io_mops_src_b; // @[Decode.scala 59:17]
  assign io_mops_write_dest = io_inst[1:0] == 2'h3 ? decoder32_io_mops_write_dest : decoder16_io_mops_write_dest; // @[Decode.scala 59:17]
  assign io_mops_alu_op = io_inst[1:0] == 2'h3 ? decoder32_io_mops_alu_op : decoder16_io_mops_alu_op; // @[Decode.scala 59:17]
  assign io_mops_alu_expand = io_inst[1:0] == 2'h3 ? decoder32_io_mops_alu_expand : decoder16_io_mops_alu_expand; // @[Decode.scala 59:17]
  assign io_mops_mem_width = io_inst[1:0] == 2'h3 ? decoder32_io_mops_mem_width : decoder16_io_mops_mem_width; // @[Decode.scala 59:17]
  assign io_mops_write_src = io_inst[1:0] == 2'h3 ? decoder32_io_mops_write_src : decoder16_io_mops_write_src; // @[Decode.scala 59:17]
  assign io_mops_rs1 = io_inst[1:0] == 2'h3 ? decoder32_io_mops_rs1 : decoder16_io_mops_rs1; // @[Decode.scala 59:17]
  assign io_mops_rs2 = io_inst[1:0] == 2'h3 ? decoder32_io_mops_rs2 : decoder16_io_mops_rs2; // @[Decode.scala 59:17]
  assign io_mops_rd = io_inst[1:0] == 2'h3 ? decoder32_io_mops_rd : decoder16_io_mops_rd; // @[Decode.scala 59:17]
  assign io_mops_imm = io_inst[1:0] == 2'h3 ? decoder32_io_mops_imm : decoder16_io_mops_imm; // @[Decode.scala 59:17]
  assign io_mops_pc = io_inst[1:0] == 2'h3 ? decoder32_io_mops_pc : decoder16_io_mops_pc; // @[Decode.scala 59:17]
  assign io_mops_predict_taken = io_inst[1:0] == 2'h3 ? decoder32_io_mops_predict_taken :
    decoder16_io_mops_predict_taken; // @[Decode.scala 59:17]
  assign io_mops_target_pc = io_inst[1:0] == 2'h3 ? decoder32_io_mops_target_pc : decoder16_io_mops_target_pc; // @[Decode.scala 59:17]
  assign io_mops_ysyx_debug = io_inst[1:0] == 2'h3 & decoder32_io_mops_ysyx_debug; // @[Decode.scala 59:17]
  assign io_mops_ysyx_print = io_inst[1:0] == 2'h3 & decoder32_io_mops_ysyx_print; // @[Decode.scala 59:17]
  assign io_mops_inst = io_inst[1:0] == 2'h3 ? decoder32_io_mops_inst : decoder16_io_mops_inst; // @[Decode.scala 59:17]
  assign decoder32_io_pc = io_pc; // @[Decode.scala 49:23]
  assign decoder32_io_inst = io_inst; // @[Decode.scala 50:23]
  assign decoder32_io_bht_predict_taken = io_bht_predict_taken; // @[Decode.scala 51:34]
  assign decoder32_io_target_pc = io_target_pc; // @[Decode.scala 52:26]
  assign decoder16_io_pc = io_pc; // @[Decode.scala 54:23]
  assign decoder16_io_inst = {{16'd0}, io_inst[15:0]}; // @[Decode.scala 55:33]
  assign decoder16_io_bht_predict_taken = io_bht_predict_taken; // @[Decode.scala 56:34]
  assign decoder16_io_target_pc = io_target_pc; // @[Decode.scala 57:26]
endmodule
module Frontend(
  input          clock,
  input          reset,
  input          io_fb_bmfs_redirect_kill,
  input  [31:0]  io_fb_bmfs_redirect_pc,
  input          io_fb_bmfs_bpu_v,
  input          io_fb_bmfs_bpu_errpr,
  input  [63:0]  io_fb_bmfs_bpu_pc_br,
  input  [63:0]  io_fb_bmfs_bpu_target,
  input          io_fb_bmfs_bpu_taken,
  output [1:0]   io_fb_fmbs_instn,
  output [160:0] io_fb_fmbs_inst_ops_0,
  output [160:0] io_fb_fmbs_inst_ops_1,
  input          io_fb_fmbs_please_wait,
  output         io_icache_req_valid,
  output [31:0]  io_icache_req_bits_addr,
  output [2:0]   io_icache_req_bits_mtype,
  input          io_icache_resp_valid,
  input  [31:0]  io_icache_resp_bits_rdata_0,
  input  [31:0]  io_icache_resp_bits_rdata_1,
  input          io_icache_resp_bits_respn,
  output         cache_stall_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  pc_gen_clock; // @[Frontend.scala 59:30]
  wire  pc_gen_reset; // @[Frontend.scala 59:30]
  wire  pc_gen_io_please_wait; // @[Frontend.scala 59:30]
  wire  pc_gen_io_redirect; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_redirect_pc; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_pc_o; // @[Frontend.scala 59:30]
  wire  pc_gen_io_predict_taken_o_0; // @[Frontend.scala 59:30]
  wire  pc_gen_io_predict_taken_o_1; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_predict_target_o_0; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_predict_target_o_1; // @[Frontend.scala 59:30]
  wire  pc_gen_io_fetch_word_o; // @[Frontend.scala 59:30]
  wire  pc_gen_io_bpu_update_dec_v; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_bpu_update_dec_pc_br; // @[Frontend.scala 59:30]
  wire  pc_gen_io_bpu_update_exe_v; // @[Frontend.scala 59:30]
  wire  pc_gen_io_bpu_update_exe_errpr; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_bpu_update_exe_pc_br; // @[Frontend.scala 59:30]
  wire [31:0] pc_gen_io_bpu_update_exe_target; // @[Frontend.scala 59:30]
  wire  pc_gen_io_bpu_update_exe_taken; // @[Frontend.scala 59:30]
  wire [31:0] Dec_io_pc; // @[Frontend.scala 70:62]
  wire [31:0] Dec_io_inst; // @[Frontend.scala 70:62]
  wire  Dec_io_bht_predict_taken; // @[Frontend.scala 70:62]
  wire [31:0] Dec_io_target_pc; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_illegal; // @[Frontend.scala 70:62]
  wire [3:0] Dec_io_mops_next_pc; // @[Frontend.scala 70:62]
  wire [1:0] Dec_io_mops_alu_mdu_lsu; // @[Frontend.scala 70:62]
  wire [3:0] Dec_io_mops_branch_type; // @[Frontend.scala 70:62]
  wire [1:0] Dec_io_mops_src_a; // @[Frontend.scala 70:62]
  wire [1:0] Dec_io_mops_src_b; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_write_dest; // @[Frontend.scala 70:62]
  wire [4:0] Dec_io_mops_alu_op; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_alu_expand; // @[Frontend.scala 70:62]
  wire [2:0] Dec_io_mops_mem_width; // @[Frontend.scala 70:62]
  wire [1:0] Dec_io_mops_write_src; // @[Frontend.scala 70:62]
  wire [4:0] Dec_io_mops_rs1; // @[Frontend.scala 70:62]
  wire [4:0] Dec_io_mops_rs2; // @[Frontend.scala 70:62]
  wire [4:0] Dec_io_mops_rd; // @[Frontend.scala 70:62]
  wire [19:0] Dec_io_mops_imm; // @[Frontend.scala 70:62]
  wire [31:0] Dec_io_mops_pc; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_predict_taken; // @[Frontend.scala 70:62]
  wire [31:0] Dec_io_mops_target_pc; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_ysyx_debug; // @[Frontend.scala 70:62]
  wire  Dec_io_mops_ysyx_print; // @[Frontend.scala 70:62]
  wire [31:0] Dec_io_mops_inst; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_pc; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_inst; // @[Frontend.scala 70:62]
  wire  Dec_1_io_bht_predict_taken; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_target_pc; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_illegal; // @[Frontend.scala 70:62]
  wire [3:0] Dec_1_io_mops_next_pc; // @[Frontend.scala 70:62]
  wire [1:0] Dec_1_io_mops_alu_mdu_lsu; // @[Frontend.scala 70:62]
  wire [3:0] Dec_1_io_mops_branch_type; // @[Frontend.scala 70:62]
  wire [1:0] Dec_1_io_mops_src_a; // @[Frontend.scala 70:62]
  wire [1:0] Dec_1_io_mops_src_b; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_write_dest; // @[Frontend.scala 70:62]
  wire [4:0] Dec_1_io_mops_alu_op; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_alu_expand; // @[Frontend.scala 70:62]
  wire [2:0] Dec_1_io_mops_mem_width; // @[Frontend.scala 70:62]
  wire [1:0] Dec_1_io_mops_write_src; // @[Frontend.scala 70:62]
  wire [4:0] Dec_1_io_mops_rs1; // @[Frontend.scala 70:62]
  wire [4:0] Dec_1_io_mops_rs2; // @[Frontend.scala 70:62]
  wire [4:0] Dec_1_io_mops_rd; // @[Frontend.scala 70:62]
  wire [19:0] Dec_1_io_mops_imm; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_mops_pc; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_predict_taken; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_mops_target_pc; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_ysyx_debug; // @[Frontend.scala 70:62]
  wire  Dec_1_io_mops_ysyx_print; // @[Frontend.scala 70:62]
  wire [31:0] Dec_1_io_mops_inst; // @[Frontend.scala 70:62]
  reg  last_req_valid; // @[Frontend.scala 61:31]
  reg [31:0] repc; // @[Frontend.scala 62:27]
  reg  renarrow; // @[Frontend.scala 63:54]
  reg [31:0] decode_pc_low_reg; // @[Frontend.scala 68:34]
  reg  decode_valid_reg; // @[Frontend.scala 69:34]
  reg  next_respn; // @[Frontend.scala 73:34]
  wire [1:0] _fire_number_respn_T = {1'h0,next_respn}; // @[Cat.scala 30:58]
  wire [1:0] fire_number_respn = _fire_number_respn_T + 2'h1; // @[Frontend.scala 74:48]
  reg [31:0] decode_pc_predict_target_0; // @[Frontend.scala 77:37]
  reg [31:0] decode_pc_predict_target_1; // @[Frontend.scala 77:37]
  reg  decode_pc_predict_taken_0; // @[Frontend.scala 78:37]
  reg  decode_pc_predict_taken_1; // @[Frontend.scala 78:37]
  reg  delayed_early_update; // @[Frontend.scala 79:37]
  wire  cache_stall = ~io_icache_resp_valid & last_req_valid; // @[Frontend.scala 92:43]
  wire  stall_f = io_fb_fmbs_please_wait | cache_stall; // @[Frontend.scala 89:29]
  reg [31:0] dec_kill_redirect_pc_REG; // @[Frontend.scala 157:34]
  wire [29:0] pc_gen_io_bpu_update_dec_pc_br_hi = decode_pc_low_reg[31:2]; // @[Frontend.scala 100:99]
  wire [1:0] pc_gen_io_bpu_update_dec_pc_br_lo = decode_pc_predict_target_0[1:0]; // @[Frontend.scala 100:145]
  wire [31:0] _pc_gen_io_bpu_update_dec_pc_br_T = {pc_gen_io_bpu_update_dec_pc_br_hi,pc_gen_io_bpu_update_dec_pc_br_lo}; // @[Cat.scala 30:58]
  wire [29:0] pc_gen_io_bpu_update_dec_pc_br_hi_1 = pc_gen_io_bpu_update_dec_pc_br_hi + 30'h1; // @[Frontend.scala 101:45]
  wire [1:0] pc_gen_io_bpu_update_dec_pc_br_lo_1 = decode_pc_predict_target_1[1:0]; // @[Frontend.scala 101:85]
  wire [31:0] _pc_gen_io_bpu_update_dec_pc_br_T_3 = {pc_gen_io_bpu_update_dec_pc_br_hi_1,
    pc_gen_io_bpu_update_dec_pc_br_lo_1}; // @[Cat.scala 30:58]
  wire  _predict_taken_but_not_br_0_T_4 = Dec_io_mops_next_pc == 4'h2 | Dec_io_mops_next_pc == 4'h3 |
    Dec_io_mops_next_pc == 4'h4; // @[Frontend.scala 83:54]
  wire  predict_taken_but_not_br_0 = Dec_io_bht_predict_taken & ~_predict_taken_but_not_br_0_T_4; // @[Frontend.scala 153:62]
  reg [31:0] pc_gen_io_bpu_update_dec_pc_br_REG; // @[Frontend.scala 100:44]
  wire [1:0] _io_icache_req_bits_mtype_T = renarrow ? 2'h2 : 2'h3; // @[Frontend.scala 124:49]
  wire [1:0] _io_icache_req_bits_mtype_T_1 = pc_gen_io_fetch_word_o ? 2'h2 : 2'h3; // @[Frontend.scala 124:89]
  wire [1:0] _io_icache_req_bits_mtype_T_2 = stall_f ? _io_icache_req_bits_mtype_T : _io_icache_req_bits_mtype_T_1; // @[Frontend.scala 124:36]
  wire  kill_d = io_fb_bmfs_redirect_kill | delayed_early_update; // @[Frontend.scala 133:39]
  wire  _GEN_5 = ~stall_f | decode_valid_reg; // @[Frontend.scala 137:25 Frontend.scala 141:30 Frontend.scala 69:34]
  wire  frontend_fire = ~cache_stall & decode_valid_reg & ~delayed_early_update; // @[Frontend.scala 144:53]
  wire [1:0] _io_fb_fmbs_instn_T_2 = decode_pc_predict_taken_0 ? 2'h1 : fire_number_respn; // @[Frontend.scala 145:62]
  wire [32:0] _T_1 = {{1'd0}, decode_pc_low_reg}; // @[Frontend.scala 148:39]
  wire [133:0] io_fb_fmbs_inst_ops_0_lo = {Dec_io_mops_rs1,Dec_io_mops_rs2,Dec_io_mops_rd,Dec_io_mops_imm,Dec_io_mops_pc
    ,Dec_io_mops_predict_taken,Dec_io_mops_target_pc,Dec_io_mops_ysyx_debug,Dec_io_mops_ysyx_print,Dec_io_mops_inst}; // @[Frontend.scala 152:44]
  wire [11:0] io_fb_fmbs_inst_ops_0_hi_lo = {Dec_io_mops_write_dest,Dec_io_mops_alu_op,Dec_io_mops_alu_expand,
    Dec_io_mops_mem_width,Dec_io_mops_write_src}; // @[Frontend.scala 152:44]
  wire [26:0] io_fb_fmbs_inst_ops_0_hi = {Dec_io_mops_illegal,Dec_io_mops_next_pc,Dec_io_mops_alu_mdu_lsu,
    Dec_io_mops_branch_type,Dec_io_mops_src_a,Dec_io_mops_src_b,io_fb_fmbs_inst_ops_0_hi_lo}; // @[Frontend.scala 152:44]
  wire [31:0] _T_4 = decode_pc_low_reg + 32'h4; // @[Frontend.scala 148:39]
  wire [133:0] io_fb_fmbs_inst_ops_1_lo = {Dec_1_io_mops_rs1,Dec_1_io_mops_rs2,Dec_1_io_mops_rd,Dec_1_io_mops_imm,
    Dec_1_io_mops_pc,Dec_1_io_mops_predict_taken,Dec_1_io_mops_target_pc,Dec_1_io_mops_ysyx_debug,
    Dec_1_io_mops_ysyx_print,Dec_1_io_mops_inst}; // @[Frontend.scala 152:44]
  wire [11:0] io_fb_fmbs_inst_ops_1_hi_lo = {Dec_1_io_mops_write_dest,Dec_1_io_mops_alu_op,Dec_1_io_mops_alu_expand,
    Dec_1_io_mops_mem_width,Dec_1_io_mops_write_src}; // @[Frontend.scala 152:44]
  wire [26:0] io_fb_fmbs_inst_ops_1_hi = {Dec_1_io_mops_illegal,Dec_1_io_mops_next_pc,Dec_1_io_mops_alu_mdu_lsu,
    Dec_1_io_mops_branch_type,Dec_1_io_mops_src_a,Dec_1_io_mops_src_b,io_fb_fmbs_inst_ops_1_hi_lo}; // @[Frontend.scala 152:44]
  wire  _predict_taken_but_not_br_1_T_4 = Dec_1_io_mops_next_pc == 4'h2 | Dec_1_io_mops_next_pc == 4'h3 |
    Dec_1_io_mops_next_pc == 4'h4; // @[Frontend.scala 83:54]
  wire  predict_taken_but_not_br_1 = Dec_1_io_bht_predict_taken & ~_predict_taken_but_not_br_1_T_4; // @[Frontend.scala 153:62]
  wire [1:0] _GEN_12 = {{1'd0}, next_respn}; // @[Frontend.scala 155:35]
  wire [1:0] _dec_update_T_2 = {predict_taken_but_not_br_1,predict_taken_but_not_br_0}; // @[Frontend.scala 155:139]
  wire  _dec_update_T_4 = _GEN_12 == 2'h0 | decode_pc_predict_taken_0 ? predict_taken_but_not_br_0 : |_dec_update_T_2; // @[Frontend.scala 155:23]
  wire  dec_update = _dec_update_T_4 & frontend_fire; // @[Frontend.scala 155:149]
  wire [31:0] _dec_kill_redirect_pc_T_3 = decode_pc_low_reg + 32'h8; // @[Frontend.scala 157:143]
  PCGen pc_gen ( // @[Frontend.scala 59:30]
    .clock(pc_gen_clock),
    .reset(pc_gen_reset),
    .io_please_wait(pc_gen_io_please_wait),
    .io_redirect(pc_gen_io_redirect),
    .io_redirect_pc(pc_gen_io_redirect_pc),
    .io_pc_o(pc_gen_io_pc_o),
    .io_predict_taken_o_0(pc_gen_io_predict_taken_o_0),
    .io_predict_taken_o_1(pc_gen_io_predict_taken_o_1),
    .io_predict_target_o_0(pc_gen_io_predict_target_o_0),
    .io_predict_target_o_1(pc_gen_io_predict_target_o_1),
    .io_fetch_word_o(pc_gen_io_fetch_word_o),
    .io_bpu_update_dec_v(pc_gen_io_bpu_update_dec_v),
    .io_bpu_update_dec_pc_br(pc_gen_io_bpu_update_dec_pc_br),
    .io_bpu_update_exe_v(pc_gen_io_bpu_update_exe_v),
    .io_bpu_update_exe_errpr(pc_gen_io_bpu_update_exe_errpr),
    .io_bpu_update_exe_pc_br(pc_gen_io_bpu_update_exe_pc_br),
    .io_bpu_update_exe_target(pc_gen_io_bpu_update_exe_target),
    .io_bpu_update_exe_taken(pc_gen_io_bpu_update_exe_taken)
  );
  Dec Dec ( // @[Frontend.scala 70:62]
    .io_pc(Dec_io_pc),
    .io_inst(Dec_io_inst),
    .io_bht_predict_taken(Dec_io_bht_predict_taken),
    .io_target_pc(Dec_io_target_pc),
    .io_mops_illegal(Dec_io_mops_illegal),
    .io_mops_next_pc(Dec_io_mops_next_pc),
    .io_mops_alu_mdu_lsu(Dec_io_mops_alu_mdu_lsu),
    .io_mops_branch_type(Dec_io_mops_branch_type),
    .io_mops_src_a(Dec_io_mops_src_a),
    .io_mops_src_b(Dec_io_mops_src_b),
    .io_mops_write_dest(Dec_io_mops_write_dest),
    .io_mops_alu_op(Dec_io_mops_alu_op),
    .io_mops_alu_expand(Dec_io_mops_alu_expand),
    .io_mops_mem_width(Dec_io_mops_mem_width),
    .io_mops_write_src(Dec_io_mops_write_src),
    .io_mops_rs1(Dec_io_mops_rs1),
    .io_mops_rs2(Dec_io_mops_rs2),
    .io_mops_rd(Dec_io_mops_rd),
    .io_mops_imm(Dec_io_mops_imm),
    .io_mops_pc(Dec_io_mops_pc),
    .io_mops_predict_taken(Dec_io_mops_predict_taken),
    .io_mops_target_pc(Dec_io_mops_target_pc),
    .io_mops_ysyx_debug(Dec_io_mops_ysyx_debug),
    .io_mops_ysyx_print(Dec_io_mops_ysyx_print),
    .io_mops_inst(Dec_io_mops_inst)
  );
  Dec Dec_1 ( // @[Frontend.scala 70:62]
    .io_pc(Dec_1_io_pc),
    .io_inst(Dec_1_io_inst),
    .io_bht_predict_taken(Dec_1_io_bht_predict_taken),
    .io_target_pc(Dec_1_io_target_pc),
    .io_mops_illegal(Dec_1_io_mops_illegal),
    .io_mops_next_pc(Dec_1_io_mops_next_pc),
    .io_mops_alu_mdu_lsu(Dec_1_io_mops_alu_mdu_lsu),
    .io_mops_branch_type(Dec_1_io_mops_branch_type),
    .io_mops_src_a(Dec_1_io_mops_src_a),
    .io_mops_src_b(Dec_1_io_mops_src_b),
    .io_mops_write_dest(Dec_1_io_mops_write_dest),
    .io_mops_alu_op(Dec_1_io_mops_alu_op),
    .io_mops_alu_expand(Dec_1_io_mops_alu_expand),
    .io_mops_mem_width(Dec_1_io_mops_mem_width),
    .io_mops_write_src(Dec_1_io_mops_write_src),
    .io_mops_rs1(Dec_1_io_mops_rs1),
    .io_mops_rs2(Dec_1_io_mops_rs2),
    .io_mops_rd(Dec_1_io_mops_rd),
    .io_mops_imm(Dec_1_io_mops_imm),
    .io_mops_pc(Dec_1_io_mops_pc),
    .io_mops_predict_taken(Dec_1_io_mops_predict_taken),
    .io_mops_target_pc(Dec_1_io_mops_target_pc),
    .io_mops_ysyx_debug(Dec_1_io_mops_ysyx_debug),
    .io_mops_ysyx_print(Dec_1_io_mops_ysyx_print),
    .io_mops_inst(Dec_1_io_mops_inst)
  );
  assign io_fb_fmbs_instn = io_fb_fmbs_please_wait | ~frontend_fire ? 2'h0 : _io_fb_fmbs_instn_T_2; // @[Frontend.scala 145:26]
  assign io_fb_fmbs_inst_ops_0 = {io_fb_fmbs_inst_ops_0_hi,io_fb_fmbs_inst_ops_0_lo}; // @[Frontend.scala 152:44]
  assign io_fb_fmbs_inst_ops_1 = {io_fb_fmbs_inst_ops_1_hi,io_fb_fmbs_inst_ops_1_lo}; // @[Frontend.scala 152:44]
  assign io_icache_req_valid = 1'h1; // @[Frontend.scala 116:28]
  assign io_icache_req_bits_addr = stall_f ? repc : pc_gen_io_pc_o; // @[Frontend.scala 118:34]
  assign io_icache_req_bits_mtype = {{1'd0}, _io_icache_req_bits_mtype_T_2}; // @[Frontend.scala 124:36]
  assign cache_stall_0 = cache_stall;
  assign pc_gen_clock = clock;
  assign pc_gen_reset = reset;
  assign pc_gen_io_please_wait = io_fb_fmbs_please_wait | cache_stall; // @[Frontend.scala 89:29]
  assign pc_gen_io_redirect = io_fb_bmfs_redirect_kill | delayed_early_update; // @[Frontend.scala 133:39]
  assign pc_gen_io_redirect_pc = io_fb_bmfs_redirect_kill ? io_fb_bmfs_redirect_pc : dec_kill_redirect_pc_REG; // @[Frontend.scala 98:31]
  assign pc_gen_io_bpu_update_dec_v = delayed_early_update; // @[Frontend.scala 102:30]
  assign pc_gen_io_bpu_update_dec_pc_br = pc_gen_io_bpu_update_dec_pc_br_REG; // @[Frontend.scala 100:34]
  assign pc_gen_io_bpu_update_exe_v = io_fb_bmfs_bpu_v; // @[Frontend.scala 103:28]
  assign pc_gen_io_bpu_update_exe_errpr = io_fb_bmfs_bpu_errpr; // @[Frontend.scala 103:28]
  assign pc_gen_io_bpu_update_exe_pc_br = io_fb_bmfs_bpu_pc_br[31:0]; // @[Frontend.scala 103:28]
  assign pc_gen_io_bpu_update_exe_target = io_fb_bmfs_bpu_target[31:0]; // @[Frontend.scala 103:28]
  assign pc_gen_io_bpu_update_exe_taken = io_fb_bmfs_bpu_taken; // @[Frontend.scala 103:28]
  assign Dec_io_pc = _T_1[31:0]; // @[Frontend.scala 148:39]
  assign Dec_io_inst = io_icache_resp_bits_rdata_0; // @[Frontend.scala 149:18]
  assign Dec_io_bht_predict_taken = decode_pc_predict_taken_0; // @[Frontend.scala 150:31]
  assign Dec_io_target_pc = decode_pc_predict_target_0; // @[Frontend.scala 151:23]
  assign Dec_1_io_pc = decode_pc_low_reg + 32'h4; // @[Frontend.scala 148:39]
  assign Dec_1_io_inst = io_icache_resp_bits_rdata_1; // @[Frontend.scala 149:18]
  assign Dec_1_io_bht_predict_taken = decode_pc_predict_taken_1; // @[Frontend.scala 150:31]
  assign Dec_1_io_target_pc = decode_pc_predict_target_1; // @[Frontend.scala 151:23]
  always @(posedge clock) begin
    if (reset) begin // @[Frontend.scala 61:31]
      last_req_valid <= 1'h0; // @[Frontend.scala 61:31]
    end else begin
      last_req_valid <= io_icache_req_valid; // @[Frontend.scala 93:18]
    end
    if (!(stall_f)) begin // @[Frontend.scala 105:14]
      repc <= pc_gen_io_pc_o;
    end
    if (!(stall_f)) begin // @[Frontend.scala 107:20]
      renarrow <= pc_gen_io_fetch_word_o;
    end
    if (reset) begin // @[Frontend.scala 68:34]
      decode_pc_low_reg <= 32'h80000000; // @[Frontend.scala 68:34]
    end else if (!(kill_d)) begin // @[Frontend.scala 135:17]
      if (~stall_f) begin // @[Frontend.scala 137:25]
        decode_pc_low_reg <= io_icache_req_bits_addr; // @[Frontend.scala 138:30]
      end
    end
    if (reset) begin // @[Frontend.scala 69:34]
      decode_valid_reg <= 1'h0; // @[Frontend.scala 69:34]
    end else if (kill_d) begin // @[Frontend.scala 135:17]
      decode_valid_reg <= 1'h0; // @[Frontend.scala 136:23]
    end else begin
      decode_valid_reg <= _GEN_5;
    end
    next_respn <= io_icache_resp_bits_respn; // @[Frontend.scala 73:34]
    if (!(kill_d)) begin // @[Frontend.scala 135:17]
      if (~stall_f) begin // @[Frontend.scala 137:25]
        decode_pc_predict_target_0 <= pc_gen_io_predict_target_o_0; // @[Frontend.scala 139:30]
      end
    end
    if (!(kill_d)) begin // @[Frontend.scala 135:17]
      if (~stall_f) begin // @[Frontend.scala 137:25]
        decode_pc_predict_target_1 <= pc_gen_io_predict_target_o_1; // @[Frontend.scala 139:30]
      end
    end
    if (!(kill_d)) begin // @[Frontend.scala 135:17]
      if (~stall_f) begin // @[Frontend.scala 137:25]
        decode_pc_predict_taken_0 <= pc_gen_io_predict_taken_o_0; // @[Frontend.scala 140:30]
      end
    end
    if (!(kill_d)) begin // @[Frontend.scala 135:17]
      if (~stall_f) begin // @[Frontend.scala 137:25]
        decode_pc_predict_taken_1 <= pc_gen_io_predict_taken_o_1; // @[Frontend.scala 140:30]
      end
    end
    if (reset) begin // @[Frontend.scala 79:37]
      delayed_early_update <= 1'h0; // @[Frontend.scala 79:37]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Frontend.scala 156:30]
      delayed_early_update <= 1'h0;
    end else begin
      delayed_early_update <= dec_update;
    end
    if (io_fb_fmbs_please_wait) begin // @[Frontend.scala 157:38]
      dec_kill_redirect_pc_REG <= decode_pc_low_reg;
    end else if (predict_taken_but_not_br_0) begin // @[Frontend.scala 157:70]
      dec_kill_redirect_pc_REG <= _T_4;
    end else begin
      dec_kill_redirect_pc_REG <= _dec_kill_redirect_pc_T_3;
    end
    if (predict_taken_but_not_br_0) begin // @[Frontend.scala 100:48]
      pc_gen_io_bpu_update_dec_pc_br_REG <= _pc_gen_io_bpu_update_dec_pc_br_T;
    end else begin
      pc_gen_io_bpu_update_dec_pc_br_REG <= _pc_gen_io_bpu_update_dec_pc_br_T_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_req_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  repc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  renarrow = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  decode_pc_low_reg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  decode_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  next_respn = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  decode_pc_predict_target_0 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  decode_pc_predict_target_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  decode_pc_predict_taken_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  decode_pc_predict_taken_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  delayed_early_update = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dec_kill_redirect_pc_REG = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  pc_gen_io_bpu_update_dec_pc_br_REG = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [63:0] io_a,
  input  [63:0] io_b,
  input  [4:0]  io_aluOp,
  input         io_aluExpand,
  input         io_aluCsr,
  input  [63:0] io_csr,
  output [63:0] io_r,
  output        io_zero
);
  wire [63:0] addResult = io_a + io_b; // @[ALU.scala 37:25]
  wire [63:0] subResult = io_a - io_b; // @[ALU.scala 38:25]
  wire [62:0] _GEN_0 = {{31'd0}, io_a[31:0]}; // @[ALU.scala 40:33]
  wire [62:0] _sllwResult_T_2 = _GEN_0 << io_b[4:0]; // @[ALU.scala 40:33]
  wire [31:0] sllwResult = _sllwResult_T_2[31:0]; // @[ALU.scala 40:47]
  wire [31:0] srlwResult = io_a[31:0] >> io_b[4:0]; // @[ALU.scala 41:32]
  wire  _T_2 = $signed(io_a) < $signed(io_b); // @[ALU.scala 45:48]
  wire  _T_4 = io_a < io_b; // @[ALU.scala 46:39]
  wire [63:0] _T_6 = io_a ^ io_b; // @[ALU.scala 47:36]
  wire [63:0] _T_7 = io_a & io_b; // @[ALU.scala 48:36]
  wire [63:0] _T_8 = io_a | io_b; // @[ALU.scala 49:36]
  wire [31:0] hi = sllwResult[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_12 = {hi,sllwResult}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_1 = {{63'd0}, io_a}; // @[ALU.scala 50:105]
  wire [126:0] _T_14 = _GEN_1 << io_b[5:0]; // @[ALU.scala 50:105]
  wire [126:0] _T_15 = io_aluExpand ? {{63'd0}, _T_12} : _T_14; // @[ALU.scala 50:33]
  wire [31:0] hi_1 = srlwResult[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_19 = {hi_1,srlwResult}; // @[Cat.scala 30:58]
  wire [63:0] _T_21 = io_a >> io_b[5:0]; // @[ALU.scala 51:105]
  wire [63:0] _T_22 = io_aluExpand ? _T_19 : _T_21; // @[ALU.scala 51:33]
  wire [31:0] hi_2 = io_a[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_27 = io_a[31:0]; // @[ALU.scala 52:100]
  wire [31:0] lo = $signed(_T_27) >>> io_b[4:0]; // @[Cat.scala 30:58]
  wire [63:0] _T_30 = {hi_2,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_34 = $signed(io_a) >>> io_b[5:0]; // @[ALU.scala 52:165]
  wire [63:0] _T_35 = io_aluExpand ? _T_30 : _T_34; // @[ALU.scala 52:33]
  wire [63:0] _alu_result_T_2 = 4'h1 == io_aluOp[3:0] ? subResult : addResult; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_4 = 4'h2 == io_aluOp[3:0] ? {{63'd0}, _T_2} : _alu_result_T_2; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_6 = 4'h3 == io_aluOp[3:0] ? {{63'd0}, _T_4} : _alu_result_T_4; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_8 = 4'h4 == io_aluOp[3:0] ? _T_6 : _alu_result_T_6; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_10 = 4'h5 == io_aluOp[3:0] ? _T_7 : _alu_result_T_8; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_12 = 4'h6 == io_aluOp[3:0] ? _T_8 : _alu_result_T_10; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_14 = 4'h7 == io_aluOp[3:0] ? _T_15 : {{63'd0}, _alu_result_T_12}; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_16 = 4'h8 == io_aluOp[3:0] ? {{63'd0}, _T_22} : _alu_result_T_14; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_18 = 4'h9 == io_aluOp[3:0] ? {{63'd0}, _T_35} : _alu_result_T_16; // @[Mux.scala 80:57]
  wire [126:0] alu_result = 4'ha == io_aluOp[3:0] ? {{63'd0}, io_b} : _alu_result_T_18; // @[Mux.scala 80:57]
  wire [31:0] alu_expand_result_hi = alu_result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_expand_result_lo = alu_result[31:0]; // @[ALU.scala 56:94]
  wire [63:0] _alu_expand_result_T_3 = {alu_expand_result_hi,alu_expand_result_lo}; // @[Cat.scala 30:58]
  wire [126:0] alu_expand_result = io_aluExpand ? {{63'd0}, _alu_expand_result_T_3} : alu_result; // @[ALU.scala 56:30]
  wire [63:0] _T_36 = io_a | io_csr; // @[ALU.scala 60:36]
  wire [63:0] _T_37 = ~io_a; // @[ALU.scala 61:36]
  wire [63:0] _T_38 = _T_37 & io_csr; // @[ALU.scala 61:52]
  wire [63:0] _csr_result_T_2 = 4'h6 == io_aluOp[3:0] ? _T_36 : io_a; // @[Mux.scala 80:57]
  wire [63:0] csr_result = 4'hb == io_aluOp[3:0] ? _T_38 : _csr_result_T_2; // @[Mux.scala 80:57]
  wire [126:0] _io_r_T = io_aluCsr ? {{63'd0}, csr_result} : alu_expand_result; // @[ALU.scala 64:16]
  assign io_r = _io_r_T[63:0]; // @[ALU.scala 64:10]
  assign io_zero = ~(|alu_expand_result); // @[ALU.scala 68:14]
endmodule
module Divider(
  input         clock,
  input         reset,
  input         io_vi,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_vo,
  output [63:0] io_div_res,
  output [63:0] io_rem_res,
  input         io_kill
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] in1d; // @[MDU.scala 149:21]
  reg [63:0] in2d; // @[MDU.scala 150:21]
  reg [1:0] state; // @[MDU.scala 153:23]
  reg [5:0] step; // @[MDU.scala 160:26]
  reg [128:0] remr; // @[MDU.scala 162:22]
  wire  isz_6 = ~(|in1d[63:56]); // @[MDU.scala 167:19]
  wire  isz_5 = ~(|in1d[55:48]); // @[MDU.scala 167:19]
  wire  isz_4 = ~(|in1d[47:40]); // @[MDU.scala 167:19]
  wire  isz_3 = ~(|in1d[39:32]); // @[MDU.scala 167:19]
  wire  isz_2 = ~(|in1d[31:24]); // @[MDU.scala 167:19]
  wire  isz_1 = ~(|in1d[23:16]); // @[MDU.scala 167:19]
  wire  isz_0 = ~(|in1d[15:8]); // @[MDU.scala 167:19]
  wire [1:0] _num_nonz_T = isz_0 ? 2'h1 : 2'h2; // @[MDU.scala 170:90]
  wire [1:0] _num_nonz_T_1 = isz_1 ? _num_nonz_T : 2'h3; // @[MDU.scala 170:78]
  wire [2:0] _num_nonz_T_2 = isz_2 ? {{1'd0}, _num_nonz_T_1} : 3'h4; // @[MDU.scala 170:66]
  wire [2:0] _num_nonz_T_3 = isz_3 ? _num_nonz_T_2 : 3'h5; // @[MDU.scala 170:54]
  wire [2:0] _num_nonz_T_4 = isz_4 ? _num_nonz_T_3 : 3'h6; // @[MDU.scala 170:42]
  wire [2:0] _num_nonz_T_5 = isz_5 ? _num_nonz_T_4 : 3'h7; // @[MDU.scala 170:30]
  wire [3:0] num_nonz = isz_6 ? {{1'd0}, _num_nonz_T_5} : 4'h8; // @[MDU.scala 170:18]
  wire [3:0] _true_rem_T_2 = 4'h8 - num_nonz; // @[MDU.scala 174:72]
  wire [7:0] _true_rem_T_3 = 4'h8 * _true_rem_T_2; // @[MDU.scala 174:52]
  wire [7:0] _true_rem_T_5 = 8'h1 + _true_rem_T_3; // @[MDU.scala 174:46]
  wire [318:0] _GEN_9 = {{255'd0}, in1d}; // @[MDU.scala 174:38]
  wire [318:0] _true_rem_T_6 = _GEN_9 << _true_rem_T_5; // @[MDU.scala 174:38]
  wire [318:0] _true_rem_T_7 = step == 6'h0 ? _true_rem_T_6 : {{190'd0}, remr}; // @[MDU.scala 174:18]
  wire [128:0] true_rem = _true_rem_T_7[128:0]; // @[MDU.scala 173:22 MDU.scala 174:12]
  wire [129:0] _rems_T_2 = {true_rem, 1'h0}; // @[MDU.scala 176:14]
  wire [63:0] _rems_T_5 = true_rem[127:64] - in2d; // @[MDU.scala 177:41]
  wire [62:0] rems_hi_hi = _rems_T_5[62:0]; // @[MDU.scala 177:48]
  wire [63:0] rems_hi_lo = true_rem[63:0]; // @[MDU.scala 177:72]
  wire [127:0] _rems_T_6 = {rems_hi_hi,rems_hi_lo,1'h1}; // @[Cat.scala 30:58]
  wire [129:0] _rems_T_7 = true_rem[127:64] < in2d ? _rems_T_2 : {{2'd0}, _rems_T_6}; // @[MDU.scala 175:18]
  wire [7:0] _nstate_T_1 = 4'h8 * num_nonz; // @[MDU.scala 187:37]
  wire [7:0] _nstate_T_3 = _nstate_T_1 - 8'h1; // @[MDU.scala 187:48]
  wire [7:0] _GEN_10 = {{2'd0}, step}; // @[MDU.scala 187:26]
  wire [1:0] _nstate_T_5 = _GEN_10 == _nstate_T_3 ? 2'h2 : 2'h1; // @[MDU.scala 187:20]
  wire [5:0] _step_T_1 = step + 6'h1; // @[MDU.scala 188:20]
  wire [128:0] rems = _rems_T_7[128:0]; // @[MDU.scala 163:23 MDU.scala 175:12]
  reg [63:0] io_div_res_REG; // @[MDU.scala 198:24]
  reg [63:0] io_rem_res_REG; // @[MDU.scala 199:24]
  assign io_vo = state == 2'h2; // @[MDU.scala 196:23]
  assign io_div_res = io_div_res_REG; // @[MDU.scala 198:14]
  assign io_rem_res = io_rem_res_REG; // @[MDU.scala 199:14]
  always @(posedge clock) begin
    in1d <= io_in1; // @[MDU.scala 149:21]
    in2d <= io_in2; // @[MDU.scala 150:21]
    if (reset) begin // @[MDU.scala 153:23]
      state <= 2'h0; // @[MDU.scala 153:23]
    end else if (state == 2'h0) begin // @[MDU.scala 180:27]
      if (io_vi) begin // @[MDU.scala 181:18]
        state <= 2'h1;
      end else begin
        state <= 2'h0;
      end
    end else if (state == 2'h1) begin // @[MDU.scala 182:32]
      if (io_kill) begin // @[MDU.scala 183:19]
        state <= 2'h0; // @[MDU.scala 184:14]
      end else begin
        state <= _nstate_T_5; // @[MDU.scala 187:14]
      end
    end else begin
      state <= 2'h0; // @[MDU.scala 193:12]
    end
    if (reset) begin // @[MDU.scala 160:26]
      step <= 6'h0; // @[MDU.scala 160:26]
    end else if (!(state == 2'h0)) begin // @[MDU.scala 180:27]
      if (state == 2'h1) begin // @[MDU.scala 182:32]
        if (io_kill) begin // @[MDU.scala 183:19]
          step <= 6'h0; // @[MDU.scala 185:12]
        end else begin
          step <= _step_T_1; // @[MDU.scala 188:12]
        end
      end else begin
        step <= 6'h0; // @[MDU.scala 192:10]
      end
    end
    if (!(state == 2'h0)) begin // @[MDU.scala 180:27]
      if (state == 2'h1) begin // @[MDU.scala 182:32]
        if (!(io_kill)) begin // @[MDU.scala 183:19]
          remr <= rems; // @[MDU.scala 189:12]
        end
      end
    end
    io_div_res_REG <= rems[63:0]; // @[MDU.scala 198:29]
    io_rem_res_REG <= rems[128:65]; // @[MDU.scala 199:29]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  in1d = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  in2d = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  step = _RAND_3[5:0];
  _RAND_4 = {5{`RANDOM}};
  remr = _RAND_4[128:0];
  _RAND_5 = {2{`RANDOM}};
  io_div_res_REG = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  io_rem_res_REG = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU_1(
  input  [63:0] io_a,
  input  [63:0] io_b,
  input  [4:0]  io_aluOp,
  input         io_aluExpand,
  output [63:0] io_r
);
  wire [63:0] addResult = io_a + io_b; // @[ALU.scala 37:25]
  wire [63:0] subResult = io_a - io_b; // @[ALU.scala 38:25]
  wire [62:0] _GEN_0 = {{31'd0}, io_a[31:0]}; // @[ALU.scala 40:33]
  wire [62:0] _sllwResult_T_2 = _GEN_0 << io_b[4:0]; // @[ALU.scala 40:33]
  wire [31:0] sllwResult = _sllwResult_T_2[31:0]; // @[ALU.scala 40:47]
  wire [31:0] srlwResult = io_a[31:0] >> io_b[4:0]; // @[ALU.scala 41:32]
  wire  _T_2 = $signed(io_a) < $signed(io_b); // @[ALU.scala 45:48]
  wire  _T_4 = io_a < io_b; // @[ALU.scala 46:39]
  wire [63:0] _T_6 = io_a ^ io_b; // @[ALU.scala 47:36]
  wire [63:0] _T_7 = io_a & io_b; // @[ALU.scala 48:36]
  wire [63:0] _T_8 = io_a | io_b; // @[ALU.scala 49:36]
  wire [31:0] hi = sllwResult[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_12 = {hi,sllwResult}; // @[Cat.scala 30:58]
  wire [126:0] _GEN_1 = {{63'd0}, io_a}; // @[ALU.scala 50:105]
  wire [126:0] _T_14 = _GEN_1 << io_b[5:0]; // @[ALU.scala 50:105]
  wire [126:0] _T_15 = io_aluExpand ? {{63'd0}, _T_12} : _T_14; // @[ALU.scala 50:33]
  wire [31:0] hi_1 = srlwResult[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_19 = {hi_1,srlwResult}; // @[Cat.scala 30:58]
  wire [63:0] _T_21 = io_a >> io_b[5:0]; // @[ALU.scala 51:105]
  wire [63:0] _T_22 = io_aluExpand ? _T_19 : _T_21; // @[ALU.scala 51:33]
  wire [31:0] hi_2 = io_a[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_27 = io_a[31:0]; // @[ALU.scala 52:100]
  wire [31:0] lo = $signed(_T_27) >>> io_b[4:0]; // @[Cat.scala 30:58]
  wire [63:0] _T_30 = {hi_2,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_34 = $signed(io_a) >>> io_b[5:0]; // @[ALU.scala 52:165]
  wire [63:0] _T_35 = io_aluExpand ? _T_30 : _T_34; // @[ALU.scala 52:33]
  wire [63:0] _alu_result_T_2 = 4'h1 == io_aluOp[3:0] ? subResult : addResult; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_4 = 4'h2 == io_aluOp[3:0] ? {{63'd0}, _T_2} : _alu_result_T_2; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_6 = 4'h3 == io_aluOp[3:0] ? {{63'd0}, _T_4} : _alu_result_T_4; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_8 = 4'h4 == io_aluOp[3:0] ? _T_6 : _alu_result_T_6; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_10 = 4'h5 == io_aluOp[3:0] ? _T_7 : _alu_result_T_8; // @[Mux.scala 80:57]
  wire [63:0] _alu_result_T_12 = 4'h6 == io_aluOp[3:0] ? _T_8 : _alu_result_T_10; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_14 = 4'h7 == io_aluOp[3:0] ? _T_15 : {{63'd0}, _alu_result_T_12}; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_16 = 4'h8 == io_aluOp[3:0] ? {{63'd0}, _T_22} : _alu_result_T_14; // @[Mux.scala 80:57]
  wire [126:0] _alu_result_T_18 = 4'h9 == io_aluOp[3:0] ? {{63'd0}, _T_35} : _alu_result_T_16; // @[Mux.scala 80:57]
  wire [126:0] alu_result = 4'ha == io_aluOp[3:0] ? {{63'd0}, io_b} : _alu_result_T_18; // @[Mux.scala 80:57]
  wire [31:0] alu_expand_result_hi = alu_result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] alu_expand_result_lo = alu_result[31:0]; // @[ALU.scala 56:94]
  wire [63:0] _alu_expand_result_T_3 = {alu_expand_result_hi,alu_expand_result_lo}; // @[Cat.scala 30:58]
  wire [126:0] alu_expand_result = io_aluExpand ? {{63'd0}, _alu_expand_result_T_3} : alu_result; // @[ALU.scala 56:30]
  assign io_r = alu_expand_result[63:0]; // @[ALU.scala 66:10]
endmodule
module MDU(
  input         clock,
  input         reset,
  input         io_kill,
  input         io_req_valid,
  input  [4:0]  io_req_op,
  input         io_req_expand,
  input  [63:0] io_req_in1,
  input  [63:0] io_req_in2,
  output [63:0] io_resp_r,
  output        io_resp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  divider_clock; // @[MDU.scala 60:23]
  wire  divider_reset; // @[MDU.scala 60:23]
  wire  divider_io_vi; // @[MDU.scala 60:23]
  wire [63:0] divider_io_in1; // @[MDU.scala 60:23]
  wire [63:0] divider_io_in2; // @[MDU.scala 60:23]
  wire  divider_io_vo; // @[MDU.scala 60:23]
  wire [63:0] divider_io_div_res; // @[MDU.scala 60:23]
  wire [63:0] divider_io_rem_res; // @[MDU.scala 60:23]
  wire  divider_io_kill; // @[MDU.scala 60:23]
  wire [63:0] alu_io_a; // @[MDU.scala 77:23]
  wire [63:0] alu_io_b; // @[MDU.scala 77:23]
  wire [4:0] alu_io_aluOp; // @[MDU.scala 77:23]
  wire  alu_io_aluExpand; // @[MDU.scala 77:23]
  wire [63:0] alu_io_r; // @[MDU.scala 77:23]
  reg [127:0] mul_res; // @[MDU.scala 51:24]
  reg [127:0] mulu_res; // @[MDU.scala 52:25]
  wire [64:0] _mulsu_res_T_1 = {1'b0,$signed(io_req_in2)}; // @[MDU.scala 53:47]
  wire [128:0] _mulsu_res_T_2 = $signed(io_req_in1) * $signed(_mulsu_res_T_1); // @[MDU.scala 53:47]
  reg [127:0] mulsu_res; // @[MDU.scala 53:26]
  wire  mdu_op = io_req_op[4]; // @[MDU.scala 55:25]
  wire  mul_op = ~io_req_op[2]; // @[MDU.scala 56:16]
  wire  div_valid = mdu_op & ~mul_op & io_req_valid; // @[MDU.scala 58:38]
  wire  mult_valid = mdu_op & mul_op & io_req_valid; // @[MDU.scala 59:37]
  wire  zerodiv = io_req_in2 == 64'h0 & div_valid; // @[MDU.scala 61:36]
  wire  overdiv = io_req_in2 == 64'hffffffffffffffff & io_req_in1 == 64'h8000000000000000 & (io_req_op == 5'h14 |
    io_req_op == 5'h16) & div_valid; // @[MDU.scala 62:168]
  wire  specialdiv = zerodiv | overdiv; // @[MDU.scala 63:28]
  reg  last_valid; // @[MDU.scala 67:27]
  wire  unsign = io_req_op == 5'h15 | io_req_op == 5'h17; // @[MDU.scala 69:42]
  wire  _sign1_T_1 = ~unsign; // @[MDU.scala 70:43]
  wire  sign1 = io_req_in1[63] & ~unsign; // @[MDU.scala 70:40]
  wire  sign2 = io_req_in2[63] & _sign1_T_1; // @[MDU.scala 71:40]
  wire [63:0] _divider_io_in1_T_1 = ~io_req_in1; // @[MDU.scala 73:41]
  wire [63:0] _divider_io_in1_T_3 = _divider_io_in1_T_1 + 64'h1; // @[MDU.scala 73:61]
  wire [63:0] _divider_io_in2_T_1 = ~io_req_in2; // @[MDU.scala 74:41]
  wire [63:0] _divider_io_in2_T_3 = _divider_io_in2_T_1 + 64'h1; // @[MDU.scala 74:61]
  wire [63:0] _result_T_6 = 2'h1 == io_req_op[1:0] ? mul_res[127:64] : mul_res[63:0]; // @[Mux.scala 80:57]
  wire [63:0] _result_T_8 = 2'h2 == io_req_op[1:0] ? mulu_res[127:64] : _result_T_6; // @[Mux.scala 80:57]
  wire [63:0] _result_T_10 = 2'h3 == io_req_op[1:0] ? mulsu_res[127:64] : _result_T_8; // @[Mux.scala 80:57]
  wire [63:0] _result_T_14 = ~divider_io_div_res; // @[MDU.scala 118:53]
  wire [63:0] _result_T_16 = _result_T_14 + 64'h1; // @[MDU.scala 118:81]
  wire [63:0] _result_T_17 = sign1 == sign2 ? divider_io_div_res : _result_T_16; // @[MDU.scala 118:14]
  wire [63:0] _result_T_19 = ~divider_io_rem_res; // @[MDU.scala 121:70]
  wire [63:0] _result_T_21 = _result_T_19 + 64'h1; // @[MDU.scala 121:98]
  wire [63:0] _result_T_22 = ~sign1 ? divider_io_rem_res : _result_T_21; // @[MDU.scala 121:39]
  wire [63:0] _result_T_24 = 2'h1 == io_req_op[1:0] ? divider_io_div_res : _result_T_17; // @[Mux.scala 80:57]
  wire [63:0] _result_T_26 = 2'h2 == io_req_op[1:0] ? _result_T_22 : _result_T_24; // @[Mux.scala 80:57]
  wire [63:0] _result_T_28 = 2'h3 == io_req_op[1:0] ? divider_io_rem_res : _result_T_26; // @[Mux.scala 80:57]
  wire [63:0] _result_res_T_5 = 2'h2 == io_req_op[1:0] ? io_req_in1 : 64'hffffffffffffffff; // @[Mux.scala 80:57]
  wire [63:0] _result_res_T_7 = 2'h3 == io_req_op[1:0] ? io_req_in1 : _result_res_T_5; // @[Mux.scala 80:57]
  wire [63:0] _result_res_T_9 = 2'h2 == io_req_op[1:0] ? 64'h0 : io_req_in1; // @[Mux.scala 80:57]
  wire [63:0] _GEN_0 = overdiv ? _result_res_T_9 : _result_T_28; // @[MDU.scala 93:26 MDU.scala 94:11 MDU.scala 99:11]
  wire [63:0] result_res = zerodiv ? _result_res_T_7 : _GEN_0; // @[MDU.scala 86:16 MDU.scala 87:11]
  wire [63:0] _result_T_29 = mul_op ? _result_T_10 : result_res; // @[MDU.scala 107:8]
  wire [63:0] result = mdu_op ? _result_T_29 : alu_io_r; // @[MDU.scala 105:16]
  wire [31:0] io_resp_r_hi = result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_resp_r_lo = result[31:0]; // @[MDU.scala 128:76]
  wire [63:0] _io_resp_r_T_3 = {io_resp_r_hi,io_resp_r_lo}; // @[Cat.scala 30:58]
  reg  mult_resp_valid_REG; // @[MDU.scala 131:44]
  wire  mult_resp_valid = ~last_valid & mult_resp_valid_REG; // @[MDU.scala 131:34]
  wire  _io_resp_valid_T_2 = mult_valid ? mult_resp_valid : 1'h1; // @[MDU.scala 132:82]
  Divider divider ( // @[MDU.scala 60:23]
    .clock(divider_clock),
    .reset(divider_reset),
    .io_vi(divider_io_vi),
    .io_in1(divider_io_in1),
    .io_in2(divider_io_in2),
    .io_vo(divider_io_vo),
    .io_div_res(divider_io_div_res),
    .io_rem_res(divider_io_rem_res),
    .io_kill(divider_io_kill)
  );
  ALU_1 alu ( // @[MDU.scala 77:23]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_aluOp(alu_io_aluOp),
    .io_aluExpand(alu_io_aluExpand),
    .io_r(alu_io_r)
  );
  assign io_resp_r = io_req_expand ? _io_resp_r_T_3 : result; // @[MDU.scala 128:19]
  assign io_resp_valid = div_valid | specialdiv ? divider_io_vo | specialdiv : _io_resp_valid_T_2; // @[MDU.scala 132:24]
  assign divider_clock = clock;
  assign divider_reset = reset;
  assign divider_io_vi = div_valid & ~zerodiv & ~overdiv; // @[MDU.scala 72:44]
  assign divider_io_in1 = sign1 ? _divider_io_in1_T_3 : io_req_in1; // @[MDU.scala 73:25]
  assign divider_io_in2 = sign2 ? _divider_io_in2_T_3 : io_req_in2; // @[MDU.scala 74:25]
  assign divider_io_kill = io_kill; // @[MDU.scala 75:19]
  assign alu_io_a = io_req_in1; // @[MDU.scala 79:19]
  assign alu_io_b = io_req_in2; // @[MDU.scala 80:19]
  assign alu_io_aluOp = io_req_op; // @[MDU.scala 81:19]
  assign alu_io_aluExpand = io_req_expand; // @[MDU.scala 82:19]
  always @(posedge clock) begin
    mul_res <= $signed(io_req_in1) * $signed(io_req_in2); // @[MDU.scala 51:43]
    mulu_res <= io_req_in1 * io_req_in2; // @[MDU.scala 52:44]
    mulsu_res <= _mulsu_res_T_2[127:0]; // @[MDU.scala 53:47]
    if (reset) begin // @[MDU.scala 67:27]
      last_valid <= 1'h0; // @[MDU.scala 67:27]
    end else begin
      last_valid <= io_resp_valid; // @[MDU.scala 130:14]
    end
    mult_resp_valid_REG <= mdu_op & mul_op & io_req_valid; // @[MDU.scala 59:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  mul_res = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  mulu_res = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  mulsu_res = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  last_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  mult_resp_valid_REG = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FIFO(
  input         clock,
  input         reset,
  output        io_dout_0_illegal,
  output [3:0]  io_dout_0_next_pc,
  output [1:0]  io_dout_0_alu_mdu_lsu,
  output [3:0]  io_dout_0_branch_type,
  output [1:0]  io_dout_0_src_a,
  output [1:0]  io_dout_0_src_b,
  output        io_dout_0_write_dest,
  output [4:0]  io_dout_0_alu_op,
  output        io_dout_0_alu_expand,
  output [2:0]  io_dout_0_mem_width,
  output [1:0]  io_dout_0_write_src,
  output [4:0]  io_dout_0_rs1,
  output [4:0]  io_dout_0_rs2,
  output [4:0]  io_dout_0_rd,
  output [19:0] io_dout_0_imm,
  output [31:0] io_dout_0_pc,
  output        io_dout_0_predict_taken,
  output [31:0] io_dout_0_target_pc,
  output        io_dout_0_ysyx_debug,
  output        io_dout_0_ysyx_print,
  output [31:0] io_dout_0_inst,
  output        io_dout_1_illegal,
  output [3:0]  io_dout_1_next_pc,
  output [1:0]  io_dout_1_alu_mdu_lsu,
  output [3:0]  io_dout_1_branch_type,
  output [1:0]  io_dout_1_src_a,
  output [1:0]  io_dout_1_src_b,
  output        io_dout_1_write_dest,
  output [4:0]  io_dout_1_alu_op,
  output        io_dout_1_alu_expand,
  output [2:0]  io_dout_1_mem_width,
  output [1:0]  io_dout_1_write_src,
  output [4:0]  io_dout_1_rs1,
  output [4:0]  io_dout_1_rs2,
  output [4:0]  io_dout_1_rd,
  output [19:0] io_dout_1_imm,
  output [31:0] io_dout_1_pc,
  output        io_dout_1_predict_taken,
  output [31:0] io_dout_1_target_pc,
  output        io_dout_1_ysyx_debug,
  output        io_dout_1_ysyx_print,
  output [31:0] io_dout_1_inst,
  input  [3:0]  io_enqStep,
  input         io_enqReq,
  input  [3:0]  io_deqStep,
  input         io_deqReq,
  input         io_din_0_illegal,
  input  [3:0]  io_din_0_next_pc,
  input  [1:0]  io_din_0_alu_mdu_lsu,
  input  [3:0]  io_din_0_branch_type,
  input  [1:0]  io_din_0_src_a,
  input  [1:0]  io_din_0_src_b,
  input         io_din_0_write_dest,
  input  [4:0]  io_din_0_alu_op,
  input         io_din_0_alu_expand,
  input  [2:0]  io_din_0_mem_width,
  input  [1:0]  io_din_0_write_src,
  input  [4:0]  io_din_0_rs1,
  input  [4:0]  io_din_0_rs2,
  input  [4:0]  io_din_0_rd,
  input  [19:0] io_din_0_imm,
  input  [31:0] io_din_0_pc,
  input         io_din_0_predict_taken,
  input  [31:0] io_din_0_target_pc,
  input         io_din_0_ysyx_debug,
  input         io_din_0_ysyx_print,
  input  [31:0] io_din_0_inst,
  input         io_din_1_illegal,
  input  [3:0]  io_din_1_next_pc,
  input  [1:0]  io_din_1_alu_mdu_lsu,
  input  [3:0]  io_din_1_branch_type,
  input  [1:0]  io_din_1_src_a,
  input  [1:0]  io_din_1_src_b,
  input         io_din_1_write_dest,
  input  [4:0]  io_din_1_alu_op,
  input         io_din_1_alu_expand,
  input  [2:0]  io_din_1_mem_width,
  input  [1:0]  io_din_1_write_src,
  input  [4:0]  io_din_1_rs1,
  input  [4:0]  io_din_1_rs2,
  input  [4:0]  io_din_1_rd,
  input  [19:0] io_din_1_imm,
  input  [31:0] io_din_1_pc,
  input         io_din_1_predict_taken,
  input  [31:0] io_din_1_target_pc,
  input         io_din_1_ysyx_debug,
  input         io_din_1_ysyx_print,
  input  [31:0] io_din_1_inst,
  input         io_flush,
  output        io_sufficient,
  output [3:0]  io_items
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
`endif // RANDOMIZE_REG_INIT
  reg  mem_0_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_0_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_0_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_0_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_0_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_0_src_b; // @[FIFO.scala 21:16]
  reg  mem_0_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_0_alu_op; // @[FIFO.scala 21:16]
  reg  mem_0_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_0_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_0_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_0_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_0_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_0_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_0_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_0_pc; // @[FIFO.scala 21:16]
  reg  mem_0_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_0_target_pc; // @[FIFO.scala 21:16]
  reg  mem_0_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_0_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_0_inst; // @[FIFO.scala 21:16]
  reg  mem_1_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_1_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_1_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_1_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_1_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_1_src_b; // @[FIFO.scala 21:16]
  reg  mem_1_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_1_alu_op; // @[FIFO.scala 21:16]
  reg  mem_1_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_1_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_1_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_1_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_1_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_1_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_1_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_1_pc; // @[FIFO.scala 21:16]
  reg  mem_1_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_1_target_pc; // @[FIFO.scala 21:16]
  reg  mem_1_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_1_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_1_inst; // @[FIFO.scala 21:16]
  reg  mem_2_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_2_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_2_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_2_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_2_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_2_src_b; // @[FIFO.scala 21:16]
  reg  mem_2_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_2_alu_op; // @[FIFO.scala 21:16]
  reg  mem_2_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_2_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_2_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_2_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_2_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_2_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_2_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_2_pc; // @[FIFO.scala 21:16]
  reg  mem_2_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_2_target_pc; // @[FIFO.scala 21:16]
  reg  mem_2_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_2_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_2_inst; // @[FIFO.scala 21:16]
  reg  mem_3_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_3_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_3_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_3_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_3_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_3_src_b; // @[FIFO.scala 21:16]
  reg  mem_3_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_3_alu_op; // @[FIFO.scala 21:16]
  reg  mem_3_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_3_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_3_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_3_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_3_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_3_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_3_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_3_pc; // @[FIFO.scala 21:16]
  reg  mem_3_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_3_target_pc; // @[FIFO.scala 21:16]
  reg  mem_3_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_3_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_3_inst; // @[FIFO.scala 21:16]
  reg  mem_4_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_4_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_4_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_4_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_4_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_4_src_b; // @[FIFO.scala 21:16]
  reg  mem_4_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_4_alu_op; // @[FIFO.scala 21:16]
  reg  mem_4_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_4_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_4_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_4_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_4_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_4_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_4_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_4_pc; // @[FIFO.scala 21:16]
  reg  mem_4_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_4_target_pc; // @[FIFO.scala 21:16]
  reg  mem_4_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_4_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_4_inst; // @[FIFO.scala 21:16]
  reg  mem_5_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_5_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_5_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_5_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_5_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_5_src_b; // @[FIFO.scala 21:16]
  reg  mem_5_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_5_alu_op; // @[FIFO.scala 21:16]
  reg  mem_5_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_5_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_5_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_5_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_5_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_5_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_5_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_5_pc; // @[FIFO.scala 21:16]
  reg  mem_5_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_5_target_pc; // @[FIFO.scala 21:16]
  reg  mem_5_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_5_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_5_inst; // @[FIFO.scala 21:16]
  reg  mem_6_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_6_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_6_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_6_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_6_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_6_src_b; // @[FIFO.scala 21:16]
  reg  mem_6_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_6_alu_op; // @[FIFO.scala 21:16]
  reg  mem_6_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_6_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_6_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_6_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_6_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_6_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_6_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_6_pc; // @[FIFO.scala 21:16]
  reg  mem_6_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_6_target_pc; // @[FIFO.scala 21:16]
  reg  mem_6_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_6_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_6_inst; // @[FIFO.scala 21:16]
  reg  mem_7_illegal; // @[FIFO.scala 21:16]
  reg [3:0] mem_7_next_pc; // @[FIFO.scala 21:16]
  reg [1:0] mem_7_alu_mdu_lsu; // @[FIFO.scala 21:16]
  reg [3:0] mem_7_branch_type; // @[FIFO.scala 21:16]
  reg [1:0] mem_7_src_a; // @[FIFO.scala 21:16]
  reg [1:0] mem_7_src_b; // @[FIFO.scala 21:16]
  reg  mem_7_write_dest; // @[FIFO.scala 21:16]
  reg [4:0] mem_7_alu_op; // @[FIFO.scala 21:16]
  reg  mem_7_alu_expand; // @[FIFO.scala 21:16]
  reg [2:0] mem_7_mem_width; // @[FIFO.scala 21:16]
  reg [1:0] mem_7_write_src; // @[FIFO.scala 21:16]
  reg [4:0] mem_7_rs1; // @[FIFO.scala 21:16]
  reg [4:0] mem_7_rs2; // @[FIFO.scala 21:16]
  reg [4:0] mem_7_rd; // @[FIFO.scala 21:16]
  reg [19:0] mem_7_imm; // @[FIFO.scala 21:16]
  reg [31:0] mem_7_pc; // @[FIFO.scala 21:16]
  reg  mem_7_predict_taken; // @[FIFO.scala 21:16]
  reg [31:0] mem_7_target_pc; // @[FIFO.scala 21:16]
  reg  mem_7_ysyx_debug; // @[FIFO.scala 21:16]
  reg  mem_7_ysyx_print; // @[FIFO.scala 21:16]
  reg [31:0] mem_7_inst; // @[FIFO.scala 21:16]
  reg  maybe_full; // @[FIFO.scala 31:27]
  reg [3:0] enqPtr; // @[FIFO.scala 24:25]
  wire [3:0] enqPtr_cntNext = enqPtr + io_enqStep; // @[FIFO.scala 25:26]
  wire [3:0] _enqPtr_cntReg_T_2 = enqPtr_cntNext - 4'h8; // @[FIFO.scala 27:48]
  wire  do_enq = io_enqReq & io_sufficient; // @[FIFO.scala 40:23]
  reg [3:0] deqPtr; // @[FIFO.scala 24:25]
  wire [3:0] deqPtr_cntNext = deqPtr + io_deqStep; // @[FIFO.scala 25:26]
  wire [3:0] _deqPtr_cntReg_T_2 = deqPtr_cntNext - 4'h8; // @[FIFO.scala 27:48]
  wire  ptr_match = enqPtr == deqPtr; // @[FIFO.scala 37:26]
  wire  empty = ptr_match & ~maybe_full | io_flush; // @[FIFO.scala 38:40]
  wire  do_deq = io_deqReq & ~empty; // @[FIFO.scala 41:23]
  wire  full = ptr_match & maybe_full; // @[FIFO.scala 39:24]
  wire [3:0] ptr_diff = enqPtr - deqPtr; // @[FIFO.scala 42:25]
  wire [3:0] _io_sufficient_T_2 = 4'h8 - io_items; // @[FIFO.scala 43:47]
  wire [3:0] _io_items_T = maybe_full ? 4'h8 : 4'h0; // @[FIFO.scala 44:33]
  wire [3:0] _io_items_T_3 = 4'h8 + ptr_diff; // @[FIFO.scala 44:88]
  wire [3:0] _io_items_T_4 = deqPtr > enqPtr ? _io_items_T_3 : ptr_diff; // @[FIFO.scala 44:63]
  wire [4:0] _T = {{1'd0}, enqPtr}; // @[FIFO.scala 48:19]
  wire [3:0] _GEN_0 = _T[3:0] % 4'h8; // @[FIFO.scala 48:26]
  wire [3:0] _T_2 = _GEN_0[3:0]; // @[FIFO.scala 48:26]
  wire [3:0] _T_5 = enqPtr + 4'h1; // @[FIFO.scala 48:19]
  wire [3:0] _GEN_1 = _T_5 % 4'h8; // @[FIFO.scala 48:26]
  wire [3:0] _T_6 = _GEN_1[3:0]; // @[FIFO.scala 48:26]
  wire [4:0] _io_dout_0_T = {{1'd0}, deqPtr}; // @[FIFO.scala 57:31]
  wire [3:0] _GEN_2 = _io_dout_0_T[3:0] % 4'h8; // @[FIFO.scala 57:38]
  wire [3:0] _io_dout_0_T_2 = _GEN_2[3:0]; // @[FIFO.scala 57:38]
  wire [31:0] _GEN_508 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_inst : mem_0_inst; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_509 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_inst : _GEN_508; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_510 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_inst : _GEN_509; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_511 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_inst : _GEN_510; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_512 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_inst : _GEN_511; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_513 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_inst : _GEN_512; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_516 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_ysyx_print : mem_0_ysyx_print; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_517 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_ysyx_print : _GEN_516; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_518 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_ysyx_print : _GEN_517; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_519 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_ysyx_print : _GEN_518; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_520 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_ysyx_print : _GEN_519; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_521 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_ysyx_print : _GEN_520; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_524 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_ysyx_debug : mem_0_ysyx_debug; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_525 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_ysyx_debug : _GEN_524; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_526 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_ysyx_debug : _GEN_525; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_527 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_ysyx_debug : _GEN_526; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_528 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_ysyx_debug : _GEN_527; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_529 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_ysyx_debug : _GEN_528; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_532 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_target_pc : mem_0_target_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_533 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_target_pc : _GEN_532; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_534 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_target_pc : _GEN_533; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_535 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_target_pc : _GEN_534; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_536 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_target_pc : _GEN_535; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_537 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_target_pc : _GEN_536; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_540 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_predict_taken : mem_0_predict_taken; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_541 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_predict_taken : _GEN_540; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_542 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_predict_taken : _GEN_541; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_543 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_predict_taken : _GEN_542; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_544 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_predict_taken : _GEN_543; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_545 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_predict_taken : _GEN_544; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_548 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_pc : mem_0_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_549 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_pc : _GEN_548; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_550 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_pc : _GEN_549; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_551 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_pc : _GEN_550; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_552 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_pc : _GEN_551; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_553 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_pc : _GEN_552; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_556 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_imm : mem_0_imm; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_557 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_imm : _GEN_556; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_558 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_imm : _GEN_557; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_559 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_imm : _GEN_558; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_560 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_imm : _GEN_559; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_561 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_imm : _GEN_560; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_564 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_rd : mem_0_rd; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_565 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_rd : _GEN_564; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_566 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_rd : _GEN_565; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_567 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_rd : _GEN_566; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_568 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_rd : _GEN_567; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_569 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_rd : _GEN_568; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_572 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_rs2 : mem_0_rs2; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_573 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_rs2 : _GEN_572; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_574 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_rs2 : _GEN_573; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_575 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_rs2 : _GEN_574; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_576 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_rs2 : _GEN_575; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_577 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_rs2 : _GEN_576; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_580 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_rs1 : mem_0_rs1; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_581 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_rs1 : _GEN_580; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_582 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_rs1 : _GEN_581; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_583 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_rs1 : _GEN_582; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_584 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_rs1 : _GEN_583; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_585 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_rs1 : _GEN_584; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_588 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_write_src : mem_0_write_src; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_589 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_write_src : _GEN_588; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_590 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_write_src : _GEN_589; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_591 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_write_src : _GEN_590; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_592 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_write_src : _GEN_591; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_593 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_write_src : _GEN_592; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_596 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_mem_width : mem_0_mem_width; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_597 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_mem_width : _GEN_596; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_598 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_mem_width : _GEN_597; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_599 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_mem_width : _GEN_598; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_600 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_mem_width : _GEN_599; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_601 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_mem_width : _GEN_600; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_604 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_alu_expand : mem_0_alu_expand; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_605 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_alu_expand : _GEN_604; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_606 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_alu_expand : _GEN_605; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_607 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_alu_expand : _GEN_606; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_608 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_alu_expand : _GEN_607; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_609 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_alu_expand : _GEN_608; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_612 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_alu_op : mem_0_alu_op; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_613 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_alu_op : _GEN_612; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_614 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_alu_op : _GEN_613; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_615 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_alu_op : _GEN_614; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_616 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_alu_op : _GEN_615; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_617 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_alu_op : _GEN_616; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_620 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_write_dest : mem_0_write_dest; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_621 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_write_dest : _GEN_620; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_622 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_write_dest : _GEN_621; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_623 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_write_dest : _GEN_622; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_624 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_write_dest : _GEN_623; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_625 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_write_dest : _GEN_624; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_628 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_src_b : mem_0_src_b; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_629 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_src_b : _GEN_628; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_630 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_src_b : _GEN_629; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_631 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_src_b : _GEN_630; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_632 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_src_b : _GEN_631; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_633 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_src_b : _GEN_632; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_636 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_src_a : mem_0_src_a; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_637 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_src_a : _GEN_636; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_638 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_src_a : _GEN_637; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_639 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_src_a : _GEN_638; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_640 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_src_a : _GEN_639; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_641 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_src_a : _GEN_640; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_644 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_branch_type : mem_0_branch_type; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_645 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_branch_type : _GEN_644; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_646 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_branch_type : _GEN_645; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_647 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_branch_type : _GEN_646; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_648 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_branch_type : _GEN_647; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_649 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_branch_type : _GEN_648; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_652 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_alu_mdu_lsu : mem_0_alu_mdu_lsu; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_653 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_alu_mdu_lsu : _GEN_652; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_654 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_alu_mdu_lsu : _GEN_653; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_655 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_alu_mdu_lsu : _GEN_654; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_656 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_alu_mdu_lsu : _GEN_655; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_657 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_alu_mdu_lsu : _GEN_656; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_660 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_next_pc : mem_0_next_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_661 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_next_pc : _GEN_660; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_662 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_next_pc : _GEN_661; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_663 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_next_pc : _GEN_662; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_664 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_next_pc : _GEN_663; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_665 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_next_pc : _GEN_664; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_668 = 3'h1 == _io_dout_0_T_2[2:0] ? mem_1_illegal : mem_0_illegal; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_669 = 3'h2 == _io_dout_0_T_2[2:0] ? mem_2_illegal : _GEN_668; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_670 = 3'h3 == _io_dout_0_T_2[2:0] ? mem_3_illegal : _GEN_669; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_671 = 3'h4 == _io_dout_0_T_2[2:0] ? mem_4_illegal : _GEN_670; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_672 = 3'h5 == _io_dout_0_T_2[2:0] ? mem_5_illegal : _GEN_671; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_673 = 3'h6 == _io_dout_0_T_2[2:0] ? mem_6_illegal : _GEN_672; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _io_dout_1_T_1 = deqPtr + 4'h1; // @[FIFO.scala 57:31]
  wire [3:0] _GEN_3 = _io_dout_1_T_1 % 4'h8; // @[FIFO.scala 57:38]
  wire [3:0] _io_dout_1_T_2 = _GEN_3[3:0]; // @[FIFO.scala 57:38]
  wire [31:0] _GEN_676 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_inst : mem_0_inst; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_677 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_inst : _GEN_676; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_678 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_inst : _GEN_677; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_679 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_inst : _GEN_678; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_680 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_inst : _GEN_679; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_681 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_inst : _GEN_680; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_684 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_ysyx_print : mem_0_ysyx_print; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_685 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_ysyx_print : _GEN_684; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_686 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_ysyx_print : _GEN_685; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_687 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_ysyx_print : _GEN_686; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_688 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_ysyx_print : _GEN_687; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_689 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_ysyx_print : _GEN_688; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_692 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_ysyx_debug : mem_0_ysyx_debug; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_693 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_ysyx_debug : _GEN_692; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_694 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_ysyx_debug : _GEN_693; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_695 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_ysyx_debug : _GEN_694; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_696 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_ysyx_debug : _GEN_695; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_697 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_ysyx_debug : _GEN_696; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_700 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_target_pc : mem_0_target_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_701 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_target_pc : _GEN_700; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_702 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_target_pc : _GEN_701; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_703 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_target_pc : _GEN_702; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_704 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_target_pc : _GEN_703; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_705 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_target_pc : _GEN_704; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_708 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_predict_taken : mem_0_predict_taken; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_709 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_predict_taken : _GEN_708; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_710 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_predict_taken : _GEN_709; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_711 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_predict_taken : _GEN_710; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_712 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_predict_taken : _GEN_711; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_713 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_predict_taken : _GEN_712; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_716 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_pc : mem_0_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_717 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_pc : _GEN_716; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_718 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_pc : _GEN_717; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_719 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_pc : _GEN_718; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_720 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_pc : _GEN_719; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [31:0] _GEN_721 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_pc : _GEN_720; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_724 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_imm : mem_0_imm; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_725 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_imm : _GEN_724; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_726 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_imm : _GEN_725; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_727 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_imm : _GEN_726; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_728 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_imm : _GEN_727; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [19:0] _GEN_729 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_imm : _GEN_728; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_732 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_rd : mem_0_rd; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_733 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_rd : _GEN_732; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_734 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_rd : _GEN_733; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_735 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_rd : _GEN_734; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_736 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_rd : _GEN_735; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_737 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_rd : _GEN_736; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_740 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_rs2 : mem_0_rs2; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_741 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_rs2 : _GEN_740; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_742 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_rs2 : _GEN_741; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_743 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_rs2 : _GEN_742; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_744 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_rs2 : _GEN_743; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_745 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_rs2 : _GEN_744; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_748 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_rs1 : mem_0_rs1; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_749 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_rs1 : _GEN_748; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_750 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_rs1 : _GEN_749; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_751 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_rs1 : _GEN_750; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_752 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_rs1 : _GEN_751; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_753 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_rs1 : _GEN_752; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_756 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_write_src : mem_0_write_src; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_757 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_write_src : _GEN_756; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_758 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_write_src : _GEN_757; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_759 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_write_src : _GEN_758; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_760 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_write_src : _GEN_759; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_761 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_write_src : _GEN_760; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_764 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_mem_width : mem_0_mem_width; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_765 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_mem_width : _GEN_764; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_766 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_mem_width : _GEN_765; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_767 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_mem_width : _GEN_766; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_768 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_mem_width : _GEN_767; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [2:0] _GEN_769 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_mem_width : _GEN_768; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_772 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_alu_expand : mem_0_alu_expand; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_773 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_alu_expand : _GEN_772; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_774 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_alu_expand : _GEN_773; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_775 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_alu_expand : _GEN_774; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_776 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_alu_expand : _GEN_775; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_777 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_alu_expand : _GEN_776; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_780 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_alu_op : mem_0_alu_op; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_781 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_alu_op : _GEN_780; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_782 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_alu_op : _GEN_781; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_783 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_alu_op : _GEN_782; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_784 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_alu_op : _GEN_783; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [4:0] _GEN_785 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_alu_op : _GEN_784; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_788 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_write_dest : mem_0_write_dest; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_789 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_write_dest : _GEN_788; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_790 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_write_dest : _GEN_789; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_791 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_write_dest : _GEN_790; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_792 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_write_dest : _GEN_791; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_793 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_write_dest : _GEN_792; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_796 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_src_b : mem_0_src_b; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_797 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_src_b : _GEN_796; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_798 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_src_b : _GEN_797; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_799 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_src_b : _GEN_798; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_800 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_src_b : _GEN_799; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_801 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_src_b : _GEN_800; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_804 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_src_a : mem_0_src_a; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_805 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_src_a : _GEN_804; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_806 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_src_a : _GEN_805; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_807 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_src_a : _GEN_806; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_808 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_src_a : _GEN_807; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_809 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_src_a : _GEN_808; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_812 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_branch_type : mem_0_branch_type; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_813 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_branch_type : _GEN_812; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_814 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_branch_type : _GEN_813; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_815 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_branch_type : _GEN_814; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_816 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_branch_type : _GEN_815; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_817 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_branch_type : _GEN_816; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_820 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_alu_mdu_lsu : mem_0_alu_mdu_lsu; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_821 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_alu_mdu_lsu : _GEN_820; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_822 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_alu_mdu_lsu : _GEN_821; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_823 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_alu_mdu_lsu : _GEN_822; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_824 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_alu_mdu_lsu : _GEN_823; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [1:0] _GEN_825 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_alu_mdu_lsu : _GEN_824; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_828 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_next_pc : mem_0_next_pc; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_829 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_next_pc : _GEN_828; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_830 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_next_pc : _GEN_829; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_831 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_next_pc : _GEN_830; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_832 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_next_pc : _GEN_831; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire [3:0] _GEN_833 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_next_pc : _GEN_832; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_836 = 3'h1 == _io_dout_1_T_2[2:0] ? mem_1_illegal : mem_0_illegal; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_837 = 3'h2 == _io_dout_1_T_2[2:0] ? mem_2_illegal : _GEN_836; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_838 = 3'h3 == _io_dout_1_T_2[2:0] ? mem_3_illegal : _GEN_837; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_839 = 3'h4 == _io_dout_1_T_2[2:0] ? mem_4_illegal : _GEN_838; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_840 = 3'h5 == _io_dout_1_T_2[2:0] ? mem_5_illegal : _GEN_839; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  wire  _GEN_841 = 3'h6 == _io_dout_1_T_2[2:0] ? mem_6_illegal : _GEN_840; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_illegal = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_illegal : _GEN_673; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_next_pc = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_next_pc : _GEN_665; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_alu_mdu_lsu = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_alu_mdu_lsu : _GEN_657; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_branch_type = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_branch_type : _GEN_649; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_src_a = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_src_a : _GEN_641; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_src_b = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_src_b : _GEN_633; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_write_dest = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_write_dest : _GEN_625; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_alu_op = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_alu_op : _GEN_617; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_alu_expand = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_alu_expand : _GEN_609; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_mem_width = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_mem_width : _GEN_601; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_write_src = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_write_src : _GEN_593; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_rs1 = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_rs1 : _GEN_585; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_rs2 = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_rs2 : _GEN_577; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_rd = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_rd : _GEN_569; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_imm = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_imm : _GEN_561; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_pc = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_pc : _GEN_553; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_predict_taken = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_predict_taken : _GEN_545; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_target_pc = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_target_pc : _GEN_537; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_ysyx_debug = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_ysyx_debug : _GEN_529; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_ysyx_print = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_ysyx_print : _GEN_521; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_0_inst = 3'h7 == _io_dout_0_T_2[2:0] ? mem_7_inst : _GEN_513; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_illegal = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_illegal : _GEN_841; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_next_pc = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_next_pc : _GEN_833; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_alu_mdu_lsu = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_alu_mdu_lsu : _GEN_825; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_branch_type = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_branch_type : _GEN_817; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_src_a = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_src_a : _GEN_809; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_src_b = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_src_b : _GEN_801; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_write_dest = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_write_dest : _GEN_793; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_alu_op = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_alu_op : _GEN_785; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_alu_expand = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_alu_expand : _GEN_777; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_mem_width = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_mem_width : _GEN_769; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_write_src = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_write_src : _GEN_761; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_rs1 = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_rs1 : _GEN_753; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_rs2 = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_rs2 : _GEN_745; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_rd = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_rd : _GEN_737; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_imm = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_imm : _GEN_729; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_pc = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_pc : _GEN_721; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_predict_taken = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_predict_taken : _GEN_713; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_target_pc = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_target_pc : _GEN_705; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_ysyx_debug = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_ysyx_debug : _GEN_697; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_ysyx_print = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_ysyx_print : _GEN_689; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_dout_1_inst = 3'h7 == _io_dout_1_T_2[2:0] ? mem_7_inst : _GEN_681; // @[FIFO.scala 57:16 FIFO.scala 57:16]
  assign io_sufficient = ~full & 4'h2 <= _io_sufficient_T_2; // @[FIFO.scala 43:26]
  assign io_items = ptr_match ? _io_items_T : _io_items_T_4; // @[FIFO.scala 44:18]
  always @(posedge clock) begin
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h0 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h0 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_0_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h1 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h1 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_1_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h2 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h2 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_2_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h3 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h3 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_3_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h4 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h4 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_4_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h5 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h5 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_5_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h6 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h6 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_6_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_illegal <= io_din_1_illegal; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_illegal <= io_din_0_illegal; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_next_pc <= io_din_1_next_pc; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_next_pc <= io_din_0_next_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_mdu_lsu <= io_din_1_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_mdu_lsu <= io_din_0_alu_mdu_lsu; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_branch_type <= io_din_1_branch_type; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_branch_type <= io_din_0_branch_type; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_src_a <= io_din_1_src_a; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_src_a <= io_din_0_src_a; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_src_b <= io_din_1_src_b; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_src_b <= io_din_0_src_b; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_write_dest <= io_din_1_write_dest; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_write_dest <= io_din_0_write_dest; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_op <= io_din_1_alu_op; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_op <= io_din_0_alu_op; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_expand <= io_din_1_alu_expand; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_alu_expand <= io_din_0_alu_expand; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_mem_width <= io_din_1_mem_width; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_mem_width <= io_din_0_mem_width; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_write_src <= io_din_1_write_src; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_write_src <= io_din_0_write_src; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rs1 <= io_din_1_rs1; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rs1 <= io_din_0_rs1; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rs2 <= io_din_1_rs2; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rs2 <= io_din_0_rs2; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rd <= io_din_1_rd; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_rd <= io_din_0_rd; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_imm <= io_din_1_imm; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_imm <= io_din_0_imm; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_pc <= io_din_1_pc; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_pc <= io_din_0_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_predict_taken <= io_din_1_predict_taken; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_predict_taken <= io_din_0_predict_taken; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_target_pc <= io_din_1_target_pc; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_target_pc <= io_din_0_target_pc; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_ysyx_debug <= io_din_1_ysyx_debug; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_ysyx_debug <= io_din_0_ysyx_debug; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_ysyx_print <= io_din_1_ysyx_print; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_ysyx_print <= io_din_0_ysyx_print; // @[FIFO.scala 48:36]
      end
    end
    if (do_enq) begin // @[FIFO.scala 46:16]
      if (3'h7 == _T_6[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_inst <= io_din_1_inst; // @[FIFO.scala 48:36]
      end else if (3'h7 == _T_2[2:0]) begin // @[FIFO.scala 48:36]
        mem_7_inst <= io_din_0_inst; // @[FIFO.scala 48:36]
      end
    end
    if (reset) begin // @[FIFO.scala 31:27]
      maybe_full <= 1'h0; // @[FIFO.scala 31:27]
    end else if (io_flush) begin // @[FIFO.scala 60:18]
      maybe_full <= 1'h0; // @[FIFO.scala 63:16]
    end else if (do_enq != do_deq) begin // @[FIFO.scala 52:27]
      maybe_full <= do_enq; // @[FIFO.scala 53:16]
    end
    if (reset) begin // @[FIFO.scala 24:25]
      enqPtr <= 4'h0; // @[FIFO.scala 24:25]
    end else if (io_flush) begin // @[FIFO.scala 60:18]
      enqPtr <= 4'h0; // @[FIFO.scala 61:12]
    end else if (do_enq) begin // @[FIFO.scala 26:16]
      if (enqPtr_cntNext >= 4'h8) begin // @[FIFO.scala 27:20]
        enqPtr <= _enqPtr_cntReg_T_2;
      end else begin
        enqPtr <= enqPtr_cntNext;
      end
    end
    if (reset) begin // @[FIFO.scala 24:25]
      deqPtr <= 4'h0; // @[FIFO.scala 24:25]
    end else if (io_flush) begin // @[FIFO.scala 60:18]
      deqPtr <= 4'h0; // @[FIFO.scala 62:12]
    end else if (do_deq) begin // @[FIFO.scala 26:16]
      if (deqPtr_cntNext >= 4'h8) begin // @[FIFO.scala 27:20]
        deqPtr <= _deqPtr_cntReg_T_2;
      end else begin
        deqPtr <= deqPtr_cntNext;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_illegal = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_next_pc = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  mem_0_alu_mdu_lsu = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  mem_0_branch_type = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  mem_0_src_a = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  mem_0_src_b = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  mem_0_write_dest = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mem_0_alu_op = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  mem_0_alu_expand = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mem_0_mem_width = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  mem_0_write_src = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  mem_0_rs1 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  mem_0_rs2 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  mem_0_rd = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  mem_0_imm = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  mem_0_pc = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_0_predict_taken = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  mem_0_target_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_0_ysyx_debug = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  mem_0_ysyx_print = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mem_0_inst = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_1_illegal = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  mem_1_next_pc = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  mem_1_alu_mdu_lsu = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  mem_1_branch_type = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  mem_1_src_a = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  mem_1_src_b = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  mem_1_write_dest = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_1_alu_op = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  mem_1_alu_expand = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mem_1_mem_width = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  mem_1_write_src = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  mem_1_rs1 = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  mem_1_rs2 = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  mem_1_rd = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  mem_1_imm = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  mem_1_pc = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mem_1_predict_taken = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  mem_1_target_pc = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mem_1_ysyx_debug = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  mem_1_ysyx_print = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  mem_1_inst = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mem_2_illegal = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  mem_2_next_pc = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  mem_2_alu_mdu_lsu = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  mem_2_branch_type = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  mem_2_src_a = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  mem_2_src_b = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  mem_2_write_dest = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  mem_2_alu_op = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  mem_2_alu_expand = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  mem_2_mem_width = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  mem_2_write_src = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  mem_2_rs1 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  mem_2_rs2 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  mem_2_rd = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  mem_2_imm = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  mem_2_pc = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  mem_2_predict_taken = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mem_2_target_pc = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mem_2_ysyx_debug = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  mem_2_ysyx_print = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  mem_2_inst = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mem_3_illegal = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  mem_3_next_pc = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  mem_3_alu_mdu_lsu = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  mem_3_branch_type = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  mem_3_src_a = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  mem_3_src_b = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  mem_3_write_dest = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  mem_3_alu_op = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  mem_3_alu_expand = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  mem_3_mem_width = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  mem_3_write_src = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  mem_3_rs1 = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  mem_3_rs2 = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  mem_3_rd = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  mem_3_imm = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  mem_3_pc = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  mem_3_predict_taken = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  mem_3_target_pc = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mem_3_ysyx_debug = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  mem_3_ysyx_print = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  mem_3_inst = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  mem_4_illegal = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  mem_4_next_pc = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  mem_4_alu_mdu_lsu = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  mem_4_branch_type = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  mem_4_src_a = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  mem_4_src_b = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  mem_4_write_dest = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  mem_4_alu_op = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  mem_4_alu_expand = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  mem_4_mem_width = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  mem_4_write_src = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  mem_4_rs1 = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  mem_4_rs2 = _RAND_96[4:0];
  _RAND_97 = {1{`RANDOM}};
  mem_4_rd = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  mem_4_imm = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  mem_4_pc = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  mem_4_predict_taken = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  mem_4_target_pc = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  mem_4_ysyx_debug = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  mem_4_ysyx_print = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  mem_4_inst = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  mem_5_illegal = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  mem_5_next_pc = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  mem_5_alu_mdu_lsu = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  mem_5_branch_type = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  mem_5_src_a = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  mem_5_src_b = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  mem_5_write_dest = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  mem_5_alu_op = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  mem_5_alu_expand = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  mem_5_mem_width = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  mem_5_write_src = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  mem_5_rs1 = _RAND_116[4:0];
  _RAND_117 = {1{`RANDOM}};
  mem_5_rs2 = _RAND_117[4:0];
  _RAND_118 = {1{`RANDOM}};
  mem_5_rd = _RAND_118[4:0];
  _RAND_119 = {1{`RANDOM}};
  mem_5_imm = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  mem_5_pc = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  mem_5_predict_taken = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  mem_5_target_pc = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  mem_5_ysyx_debug = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  mem_5_ysyx_print = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  mem_5_inst = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  mem_6_illegal = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  mem_6_next_pc = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  mem_6_alu_mdu_lsu = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  mem_6_branch_type = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  mem_6_src_a = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  mem_6_src_b = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  mem_6_write_dest = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  mem_6_alu_op = _RAND_133[4:0];
  _RAND_134 = {1{`RANDOM}};
  mem_6_alu_expand = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  mem_6_mem_width = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  mem_6_write_src = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  mem_6_rs1 = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  mem_6_rs2 = _RAND_138[4:0];
  _RAND_139 = {1{`RANDOM}};
  mem_6_rd = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  mem_6_imm = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  mem_6_pc = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  mem_6_predict_taken = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  mem_6_target_pc = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  mem_6_ysyx_debug = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  mem_6_ysyx_print = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  mem_6_inst = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  mem_7_illegal = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  mem_7_next_pc = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  mem_7_alu_mdu_lsu = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  mem_7_branch_type = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  mem_7_src_a = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  mem_7_src_b = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  mem_7_write_dest = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  mem_7_alu_op = _RAND_154[4:0];
  _RAND_155 = {1{`RANDOM}};
  mem_7_alu_expand = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  mem_7_mem_width = _RAND_156[2:0];
  _RAND_157 = {1{`RANDOM}};
  mem_7_write_src = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  mem_7_rs1 = _RAND_158[4:0];
  _RAND_159 = {1{`RANDOM}};
  mem_7_rs2 = _RAND_159[4:0];
  _RAND_160 = {1{`RANDOM}};
  mem_7_rd = _RAND_160[4:0];
  _RAND_161 = {1{`RANDOM}};
  mem_7_imm = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  mem_7_pc = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  mem_7_predict_taken = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  mem_7_target_pc = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  mem_7_ysyx_debug = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  mem_7_ysyx_print = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  mem_7_inst = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  maybe_full = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  enqPtr = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  deqPtr = _RAND_170[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IssueArbiter(
  input         io_insts_in_0_illegal,
  input  [3:0]  io_insts_in_0_next_pc,
  input  [1:0]  io_insts_in_0_alu_mdu_lsu,
  input  [3:0]  io_insts_in_0_branch_type,
  input  [1:0]  io_insts_in_0_src_a,
  input  [1:0]  io_insts_in_0_src_b,
  input         io_insts_in_0_write_dest,
  input  [4:0]  io_insts_in_0_alu_op,
  input         io_insts_in_0_alu_expand,
  input  [2:0]  io_insts_in_0_mem_width,
  input  [1:0]  io_insts_in_0_write_src,
  input  [4:0]  io_insts_in_0_rs1,
  input  [4:0]  io_insts_in_0_rs2,
  input  [4:0]  io_insts_in_0_rd,
  input  [19:0] io_insts_in_0_imm,
  input  [31:0] io_insts_in_0_pc,
  input         io_insts_in_0_predict_taken,
  input  [31:0] io_insts_in_0_target_pc,
  input         io_insts_in_0_ysyx_debug,
  input         io_insts_in_0_ysyx_print,
  input  [31:0] io_insts_in_0_inst,
  input         io_insts_in_1_illegal,
  input  [3:0]  io_insts_in_1_next_pc,
  input  [1:0]  io_insts_in_1_alu_mdu_lsu,
  input  [3:0]  io_insts_in_1_branch_type,
  input  [1:0]  io_insts_in_1_src_a,
  input  [1:0]  io_insts_in_1_src_b,
  input         io_insts_in_1_write_dest,
  input  [4:0]  io_insts_in_1_alu_op,
  input         io_insts_in_1_alu_expand,
  input  [2:0]  io_insts_in_1_mem_width,
  input  [1:0]  io_insts_in_1_write_src,
  input  [4:0]  io_insts_in_1_rs1,
  input  [4:0]  io_insts_in_1_rs2,
  input  [4:0]  io_insts_in_1_rd,
  input  [19:0] io_insts_in_1_imm,
  input  [31:0] io_insts_in_1_pc,
  input         io_insts_in_1_predict_taken,
  input  [31:0] io_insts_in_1_target_pc,
  input         io_insts_in_1_ysyx_debug,
  input         io_insts_in_1_ysyx_print,
  input  [31:0] io_insts_in_1_inst,
  input  [3:0]  io_queue_items,
  input  [4:0]  io_ld_dest_ex,
  input  [63:0] io_rss_in_0,
  input  [63:0] io_rss_in_1,
  input  [63:0] io_rts_in_0,
  input  [63:0] io_rts_in_1,
  output [63:0] io_rss_out_0,
  output [63:0] io_rss_out_1,
  output [63:0] io_rss_out_2,
  output [63:0] io_rts_out_0,
  output [63:0] io_rts_out_1,
  output [63:0] io_rts_out_2,
  output        io_insts_out_0_illegal,
  output [3:0]  io_insts_out_0_next_pc,
  output [1:0]  io_insts_out_0_alu_mdu_lsu,
  output [3:0]  io_insts_out_0_branch_type,
  output [1:0]  io_insts_out_0_src_a,
  output [1:0]  io_insts_out_0_src_b,
  output        io_insts_out_0_write_dest,
  output [4:0]  io_insts_out_0_alu_op,
  output        io_insts_out_0_alu_expand,
  output [1:0]  io_insts_out_0_write_src,
  output [4:0]  io_insts_out_0_rs1,
  output [4:0]  io_insts_out_0_rd,
  output [19:0] io_insts_out_0_imm,
  output [31:0] io_insts_out_0_pc,
  output        io_insts_out_0_predict_taken,
  output [31:0] io_insts_out_0_target_pc,
  output        io_insts_out_0_ysyx_debug,
  output        io_insts_out_0_ysyx_print,
  output [31:0] io_insts_out_0_inst,
  output [1:0]  io_insts_out_1_src_a,
  output [1:0]  io_insts_out_1_src_b,
  output        io_insts_out_1_write_dest,
  output [4:0]  io_insts_out_1_alu_op,
  output        io_insts_out_1_alu_expand,
  output [4:0]  io_insts_out_1_rd,
  output [19:0] io_insts_out_1_imm,
  output [31:0] io_insts_out_1_pc,
  output        io_insts_out_1_ysyx_print,
  output [31:0] io_insts_out_1_inst,
  output [1:0]  io_insts_out_2_src_a,
  output        io_insts_out_2_write_dest,
  output [4:0]  io_insts_out_2_alu_op,
  output [2:0]  io_insts_out_2_mem_width,
  output [4:0]  io_insts_out_2_rd,
  output [19:0] io_insts_out_2_imm,
  output [31:0] io_insts_out_2_pc,
  output        io_insts_out_2_ysyx_print,
  output [31:0] io_insts_out_2_inst,
  output [1:0]  io_issue_num,
  output        io_issue_fu_valid_0,
  output        io_issue_fu_valid_1,
  output        io_issue_fu_valid_2,
  output [1:0]  io_insts_order_0,
  output [1:0]  io_insts_order_1,
  output [1:0]  io_insts_order_2
);
  wire  _T_5 = io_ld_dest_ex == 5'h0 | io_insts_in_0_rs1 != io_ld_dest_ex & io_insts_in_0_rs2 != io_ld_dest_ex; // @[IssueArbiter.scala 39:18]
  wire  issue_valid_0 = io_queue_items > 4'h0 & _T_5; // @[IssueArbiter.scala 53:29]
  wire  _T_8 = io_insts_in_0_rd != 5'h0; // @[IssueArbiter.scala 31:14]
  wire  _T_12 = io_insts_in_0_rd != 5'h0 & (io_insts_in_0_rd == io_insts_in_1_rs1 | io_insts_in_0_rd ==
    io_insts_in_1_rs2); // @[IssueArbiter.scala 31:22]
  wire  _T_15 = _T_8 & io_insts_in_0_rd == io_insts_in_1_rd; // @[IssueArbiter.scala 27:22]
  wire  _T_16 = _T_12 | _T_15; // @[IssueArbiter.scala 35:25]
  wire  _T_19 = io_insts_in_0_alu_mdu_lsu == 2'h3; // @[IssueArbiter.scala 45:29]
  wire  _T_20 = io_insts_in_1_alu_mdu_lsu == 2'h3; // @[IssueArbiter.scala 45:62]
  wire  _T_21 = io_insts_in_0_alu_mdu_lsu == 2'h3 & io_insts_in_1_alu_mdu_lsu == 2'h3; // @[IssueArbiter.scala 45:41]
  wire  _T_22 = io_insts_in_0_alu_mdu_lsu != io_insts_in_1_alu_mdu_lsu | _T_21; // @[IssueArbiter.scala 44:48]
  wire  _T_23 = ~_T_16 & _T_22; // @[IssueArbiter.scala 43:33]
  wire  _T_33 = ~(io_insts_in_0_alu_mdu_lsu == 2'h2 & io_insts_in_1_alu_mdu_lsu == 2'h1 | io_insts_in_0_alu_mdu_lsu == 2'h1
     & io_insts_in_1_alu_mdu_lsu == 2'h2); // @[IssueArbiter.scala 46:7]
  wire  _T_34 = _T_23 & io_insts_in_0_alu_mdu_lsu != 2'h0 & _T_33; // @[IssueArbiter.scala 45:108]
  wire  _T_40 = io_ld_dest_ex == 5'h0 | io_insts_in_1_rs1 != io_ld_dest_ex & io_insts_in_1_rs2 != io_ld_dest_ex; // @[IssueArbiter.scala 39:18]
  wire  _T_41 = io_queue_items > 4'h1 & _T_34 & _T_40; // @[IssueArbiter.scala 56:79]
  wire [1:0] _GEN_1 = _T_41 ? 2'h2 : 2'h1; // @[IssueArbiter.scala 57:58 IssueArbiter.scala 60:20 IssueArbiter.scala 55:18]
  wire  issue_valid_1 = issue_valid_0 & _T_41; // @[IssueArbiter.scala 53:83]
  wire  _T_42 = 2'h0 == io_insts_in_0_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire  _T_43 = 2'h1 == io_insts_in_0_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire  _T_44 = 2'h2 == io_insts_in_0_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_5 = _T_44 ? io_insts_in_0_inst : 32'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire  _GEN_6 = _T_44 & io_insts_in_0_ysyx_print; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_10 = _T_44 ? io_insts_in_0_pc : 32'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_11 = _T_44 ? io_insts_in_0_imm : 20'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_12 = _T_44 ? io_insts_in_0_rd : 5'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [2:0] _GEN_16 = _T_44 ? io_insts_in_0_mem_width : 3'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_18 = _T_44 ? io_insts_in_0_alu_op : 5'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire  _GEN_19 = _T_44 & io_insts_in_0_write_dest; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_21 = _T_44 ? io_insts_in_0_src_a : 2'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_26 = _T_44 ? io_rss_in_0 : 64'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 98:25 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_27 = _T_44 ? io_rts_in_0 : 64'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 99:25 IssueArbiter.scala 73:19]
  wire [31:0] _GEN_30 = _T_43 ? io_insts_in_0_inst : 32'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire  _GEN_31 = _T_43 & io_insts_in_0_ysyx_print; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_35 = _T_43 ? io_insts_in_0_pc : 32'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_36 = _T_43 ? io_insts_in_0_imm : 20'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_37 = _T_43 ? io_insts_in_0_rd : 5'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire  _GEN_42 = _T_43 & io_insts_in_0_alu_expand; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_43 = _T_43 ? io_insts_in_0_alu_op : 5'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire  _GEN_44 = _T_43 & io_insts_in_0_write_dest; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_45 = _T_43 ? io_insts_in_0_src_b : 2'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_46 = _T_43 ? io_insts_in_0_src_a : 2'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_51 = _T_43 ? io_rss_in_0 : 64'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 90:25 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_52 = _T_43 ? io_rts_in_0 : 64'h0; // @[Conditional.scala 39:67 IssueArbiter.scala 91:25 IssueArbiter.scala 73:19]
  wire [31:0] _GEN_55 = _T_43 ? 32'h0 : _GEN_5; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire  _GEN_56 = _T_43 ? 1'h0 : _GEN_6; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_60 = _T_43 ? 32'h0 : _GEN_10; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_61 = _T_43 ? 20'h0 : _GEN_11; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_62 = _T_43 ? 5'h0 : _GEN_12; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [2:0] _GEN_66 = _T_43 ? 3'h0 : _GEN_16; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_68 = _T_43 ? 5'h0 : _GEN_18; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire  _GEN_69 = _T_43 ? 1'h0 : _GEN_19; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_71 = _T_43 ? 2'h0 : _GEN_21; // @[Conditional.scala 39:67 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_76 = _T_43 ? 64'h0 : _GEN_26; // @[Conditional.scala 39:67 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_77 = _T_43 ? 64'h0 : _GEN_27; // @[Conditional.scala 39:67 IssueArbiter.scala 73:19]
  wire  _GEN_79 = _T_43 ? 1'h0 : _T_44; // @[Conditional.scala 39:67 IssueArbiter.scala 75:26]
  wire [31:0] _GEN_80 = _T_42 ? io_insts_in_0_inst : 32'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_81 = _T_42 & io_insts_in_0_ysyx_print; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_82 = _T_42 & io_insts_in_0_ysyx_debug; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_83 = _T_42 ? io_insts_in_0_target_pc : 32'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_84 = _T_42 & io_insts_in_0_predict_taken; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_85 = _T_42 ? io_insts_in_0_pc : 32'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_86 = _T_42 ? io_insts_in_0_imm : 20'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_87 = _T_42 ? io_insts_in_0_rd : 5'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_89 = _T_42 ? io_insts_in_0_rs1 : 5'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_90 = _T_42 ? io_insts_in_0_write_src : 2'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_92 = _T_42 & io_insts_in_0_alu_expand; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_93 = _T_42 ? io_insts_in_0_alu_op : 5'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_94 = _T_42 & io_insts_in_0_write_dest; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_95 = _T_42 ? io_insts_in_0_src_b : 2'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_96 = _T_42 ? io_insts_in_0_src_a : 2'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [3:0] _GEN_97 = _T_42 ? io_insts_in_0_branch_type : 4'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_98 = _T_42 ? io_insts_in_0_alu_mdu_lsu : 2'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [3:0] _GEN_99 = _T_42 ? io_insts_in_0_next_pc : 4'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire  _GEN_100 = _T_42 & io_insts_in_0_illegal; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_101 = _T_42 ? io_rss_in_0 : 64'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 82:25 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_102 = _T_42 ? io_rts_in_0 : 64'h0; // @[Conditional.scala 40:58 IssueArbiter.scala 83:25 IssueArbiter.scala 73:19]
  wire [31:0] _GEN_105 = _T_42 ? 32'h0 : _GEN_30; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire  _GEN_106 = _T_42 ? 1'h0 : _GEN_31; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_110 = _T_42 ? 32'h0 : _GEN_35; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_111 = _T_42 ? 20'h0 : _GEN_36; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_112 = _T_42 ? 5'h0 : _GEN_37; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire  _GEN_117 = _T_42 ? 1'h0 : _GEN_42; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_118 = _T_42 ? 5'h0 : _GEN_43; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire  _GEN_119 = _T_42 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_120 = _T_42 ? 2'h0 : _GEN_45; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_121 = _T_42 ? 2'h0 : _GEN_46; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_126 = _T_42 ? 64'h0 : _GEN_51; // @[Conditional.scala 40:58 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_127 = _T_42 ? 64'h0 : _GEN_52; // @[Conditional.scala 40:58 IssueArbiter.scala 73:19]
  wire  _GEN_129 = _T_42 ? 1'h0 : _T_43; // @[Conditional.scala 40:58 IssueArbiter.scala 75:26]
  wire [31:0] _GEN_130 = _T_42 ? 32'h0 : _GEN_55; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire  _GEN_131 = _T_42 ? 1'h0 : _GEN_56; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_135 = _T_42 ? 32'h0 : _GEN_60; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_136 = _T_42 ? 20'h0 : _GEN_61; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_137 = _T_42 ? 5'h0 : _GEN_62; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [2:0] _GEN_141 = _T_42 ? 3'h0 : _GEN_66; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_143 = _T_42 ? 5'h0 : _GEN_68; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire  _GEN_144 = _T_42 ? 1'h0 : _GEN_69; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_146 = _T_42 ? 2'h0 : _GEN_71; // @[Conditional.scala 40:58 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_151 = _T_42 ? 64'h0 : _GEN_76; // @[Conditional.scala 40:58 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_152 = _T_42 ? 64'h0 : _GEN_77; // @[Conditional.scala 40:58 IssueArbiter.scala 73:19]
  wire  _GEN_154 = _T_42 ? 1'h0 : _GEN_79; // @[Conditional.scala 40:58 IssueArbiter.scala 75:26]
  wire [31:0] _GEN_155 = issue_valid_0 ? _GEN_80 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_156 = issue_valid_0 & _GEN_81; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_157 = issue_valid_0 & _GEN_82; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_158 = issue_valid_0 ? _GEN_83 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_159 = issue_valid_0 & _GEN_84; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_160 = issue_valid_0 ? _GEN_85 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_161 = issue_valid_0 ? _GEN_86 : 20'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_162 = issue_valid_0 ? _GEN_87 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_164 = issue_valid_0 ? _GEN_89 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_165 = issue_valid_0 ? _GEN_90 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_167 = issue_valid_0 & _GEN_92; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_168 = issue_valid_0 ? _GEN_93 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_169 = issue_valid_0 & _GEN_94; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_170 = issue_valid_0 ? _GEN_95 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_171 = issue_valid_0 ? _GEN_96 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [3:0] _GEN_172 = issue_valid_0 ? _GEN_97 : 4'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_173 = issue_valid_0 ? _GEN_98 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [3:0] _GEN_174 = issue_valid_0 ? _GEN_99 : 4'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_175 = issue_valid_0 & _GEN_100; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_176 = issue_valid_0 ? _GEN_101 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_177 = issue_valid_0 ? _GEN_102 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 73:19]
  wire  _GEN_179 = issue_valid_0 & _T_42; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 75:26]
  wire [31:0] _GEN_180 = issue_valid_0 ? _GEN_105 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_181 = issue_valid_0 & _GEN_106; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_185 = issue_valid_0 ? _GEN_110 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_186 = issue_valid_0 ? _GEN_111 : 20'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_187 = issue_valid_0 ? _GEN_112 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_192 = issue_valid_0 & _GEN_117; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_193 = issue_valid_0 ? _GEN_118 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_194 = issue_valid_0 & _GEN_119; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_195 = issue_valid_0 ? _GEN_120 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_196 = issue_valid_0 ? _GEN_121 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_201 = issue_valid_0 ? _GEN_126 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_202 = issue_valid_0 ? _GEN_127 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 73:19]
  wire  _GEN_204 = issue_valid_0 & _GEN_129; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 75:26]
  wire [31:0] _GEN_205 = issue_valid_0 ? _GEN_130 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_206 = issue_valid_0 & _GEN_131; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [31:0] _GEN_210 = issue_valid_0 ? _GEN_135 : 32'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [19:0] _GEN_211 = issue_valid_0 ? _GEN_136 : 20'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_212 = issue_valid_0 ? _GEN_137 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [2:0] _GEN_216 = issue_valid_0 ? _GEN_141 : 3'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [4:0] _GEN_218 = issue_valid_0 ? _GEN_143 : 5'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire  _GEN_219 = issue_valid_0 & _GEN_144; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [1:0] _GEN_221 = issue_valid_0 ? _GEN_146 : 2'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 71:21]
  wire [63:0] _GEN_226 = issue_valid_0 ? _GEN_151 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 72:19]
  wire [63:0] _GEN_227 = issue_valid_0 ? _GEN_152 : 64'h0; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 73:19]
  wire  _GEN_229 = issue_valid_0 & _GEN_154; // @[IssueArbiter.scala 78:26 IssueArbiter.scala 75:26]
  wire  _T_53 = 2'h0 == io_insts_in_1_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire  _GEN_581 = _T_53 | _GEN_179; // @[Conditional.scala 40:58 IssueArbiter.scala 86:22]
  wire  alu_occupy = issue_valid_1 ? _GEN_581 : _GEN_179; // @[IssueArbiter.scala 78:26]
  wire  _T_47 = ~alu_occupy; // @[IssueArbiter.scala 108:14]
  wire  _T_54 = 2'h1 == io_insts_in_1_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire  _GEN_530 = _T_54 | _GEN_204; // @[Conditional.scala 39:67 IssueArbiter.scala 94:22]
  wire  _GEN_607 = _T_53 ? _GEN_204 : _GEN_530; // @[Conditional.scala 40:58]
  wire  mdu_occupy = issue_valid_1 ? _GEN_607 : _GEN_204; // @[IssueArbiter.scala 78:26]
  wire  _T_48 = ~mdu_occupy; // @[IssueArbiter.scala 114:21]
  wire [31:0] _GEN_230 = ~mdu_occupy ? io_insts_in_0_inst : _GEN_180; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_231 = ~mdu_occupy ? io_insts_in_0_ysyx_print : _GEN_181; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [31:0] _GEN_235 = ~mdu_occupy ? io_insts_in_0_pc : _GEN_185; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [19:0] _GEN_236 = ~mdu_occupy ? io_insts_in_0_imm : _GEN_186; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_237 = ~mdu_occupy ? io_insts_in_0_rd : _GEN_187; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_242 = ~mdu_occupy ? io_insts_in_0_alu_expand : _GEN_192; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_243 = ~mdu_occupy ? io_insts_in_0_alu_op : _GEN_193; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_244 = ~mdu_occupy ? io_insts_in_0_write_dest : _GEN_194; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_245 = ~mdu_occupy ? io_insts_in_0_src_b : _GEN_195; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_246 = ~mdu_occupy ? io_insts_in_0_src_a : _GEN_196; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [63:0] _GEN_251 = ~mdu_occupy ? io_rss_in_0 : _GEN_201; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 116:25]
  wire [63:0] _GEN_252 = ~mdu_occupy ? io_rts_in_0 : _GEN_202; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 117:25]
  wire  _GEN_254 = ~mdu_occupy | _GEN_204; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 119:32]
  wire [31:0] _GEN_255 = ~alu_occupy ? io_insts_in_0_inst : _GEN_155; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_256 = ~alu_occupy ? io_insts_in_0_ysyx_print : _GEN_156; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_257 = ~alu_occupy ? io_insts_in_0_ysyx_debug : _GEN_157; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_258 = ~alu_occupy ? io_insts_in_0_target_pc : _GEN_158; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_259 = ~alu_occupy ? io_insts_in_0_predict_taken : _GEN_159; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_260 = ~alu_occupy ? io_insts_in_0_pc : _GEN_160; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [19:0] _GEN_261 = ~alu_occupy ? io_insts_in_0_imm : _GEN_161; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_262 = ~alu_occupy ? io_insts_in_0_rd : _GEN_162; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_264 = ~alu_occupy ? io_insts_in_0_rs1 : _GEN_164; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_265 = ~alu_occupy ? io_insts_in_0_write_src : _GEN_165; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_267 = ~alu_occupy ? io_insts_in_0_alu_expand : _GEN_167; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_268 = ~alu_occupy ? io_insts_in_0_alu_op : _GEN_168; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_269 = ~alu_occupy ? io_insts_in_0_write_dest : _GEN_169; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_270 = ~alu_occupy ? io_insts_in_0_src_b : _GEN_170; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_271 = ~alu_occupy ? io_insts_in_0_src_a : _GEN_171; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_272 = ~alu_occupy ? io_insts_in_0_branch_type : _GEN_172; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_273 = ~alu_occupy ? io_insts_in_0_alu_mdu_lsu : _GEN_173; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_274 = ~alu_occupy ? io_insts_in_0_next_pc : _GEN_174; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_275 = ~alu_occupy ? io_insts_in_0_illegal : _GEN_175; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [63:0] _GEN_276 = ~alu_occupy ? io_rss_in_0 : _GEN_176; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 110:25]
  wire [63:0] _GEN_277 = ~alu_occupy ? io_rts_in_0 : _GEN_177; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 111:25]
  wire  _GEN_279 = ~alu_occupy | _GEN_179; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 113:32]
  wire [31:0] _GEN_280 = ~alu_occupy ? _GEN_180 : _GEN_230; // @[IssueArbiter.scala 108:27]
  wire  _GEN_281 = ~alu_occupy ? _GEN_181 : _GEN_231; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_285 = ~alu_occupy ? _GEN_185 : _GEN_235; // @[IssueArbiter.scala 108:27]
  wire [19:0] _GEN_286 = ~alu_occupy ? _GEN_186 : _GEN_236; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_287 = ~alu_occupy ? _GEN_187 : _GEN_237; // @[IssueArbiter.scala 108:27]
  wire  _GEN_292 = ~alu_occupy ? _GEN_192 : _GEN_242; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_293 = ~alu_occupy ? _GEN_193 : _GEN_243; // @[IssueArbiter.scala 108:27]
  wire  _GEN_294 = ~alu_occupy ? _GEN_194 : _GEN_244; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_295 = ~alu_occupy ? _GEN_195 : _GEN_245; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_296 = ~alu_occupy ? _GEN_196 : _GEN_246; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_301 = ~alu_occupy ? _GEN_201 : _GEN_251; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_302 = ~alu_occupy ? _GEN_202 : _GEN_252; // @[IssueArbiter.scala 108:27]
  wire  _GEN_304 = ~alu_occupy ? _GEN_204 : _GEN_254; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_305 = issue_valid_0 & _T_19 ? _GEN_255 : _GEN_155; // @[IssueArbiter.scala 107:70]
  wire  _GEN_306 = issue_valid_0 & _T_19 ? _GEN_256 : _GEN_156; // @[IssueArbiter.scala 107:70]
  wire  _GEN_307 = issue_valid_0 & _T_19 ? _GEN_257 : _GEN_157; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_308 = issue_valid_0 & _T_19 ? _GEN_258 : _GEN_158; // @[IssueArbiter.scala 107:70]
  wire  _GEN_309 = issue_valid_0 & _T_19 ? _GEN_259 : _GEN_159; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_310 = issue_valid_0 & _T_19 ? _GEN_260 : _GEN_160; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_311 = issue_valid_0 & _T_19 ? _GEN_261 : _GEN_161; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_312 = issue_valid_0 & _T_19 ? _GEN_262 : _GEN_162; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_314 = issue_valid_0 & _T_19 ? _GEN_264 : _GEN_164; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_315 = issue_valid_0 & _T_19 ? _GEN_265 : _GEN_165; // @[IssueArbiter.scala 107:70]
  wire  _GEN_317 = issue_valid_0 & _T_19 ? _GEN_267 : _GEN_167; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_318 = issue_valid_0 & _T_19 ? _GEN_268 : _GEN_168; // @[IssueArbiter.scala 107:70]
  wire  _GEN_319 = issue_valid_0 & _T_19 ? _GEN_269 : _GEN_169; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_320 = issue_valid_0 & _T_19 ? _GEN_270 : _GEN_170; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_321 = issue_valid_0 & _T_19 ? _GEN_271 : _GEN_171; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_322 = issue_valid_0 & _T_19 ? _GEN_272 : _GEN_172; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_323 = issue_valid_0 & _T_19 ? _GEN_273 : _GEN_173; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_324 = issue_valid_0 & _T_19 ? _GEN_274 : _GEN_174; // @[IssueArbiter.scala 107:70]
  wire  _GEN_325 = issue_valid_0 & _T_19 ? _GEN_275 : _GEN_175; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_326 = issue_valid_0 & _T_19 ? _GEN_276 : _GEN_176; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_327 = issue_valid_0 & _T_19 ? _GEN_277 : _GEN_177; // @[IssueArbiter.scala 107:70]
  wire  _GEN_329 = issue_valid_0 & _T_19 ? _GEN_279 : _GEN_179; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_330 = issue_valid_0 & _T_19 ? _GEN_280 : _GEN_180; // @[IssueArbiter.scala 107:70]
  wire  _GEN_331 = issue_valid_0 & _T_19 ? _GEN_281 : _GEN_181; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_335 = issue_valid_0 & _T_19 ? _GEN_285 : _GEN_185; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_336 = issue_valid_0 & _T_19 ? _GEN_286 : _GEN_186; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_337 = issue_valid_0 & _T_19 ? _GEN_287 : _GEN_187; // @[IssueArbiter.scala 107:70]
  wire  _GEN_342 = issue_valid_0 & _T_19 ? _GEN_292 : _GEN_192; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_343 = issue_valid_0 & _T_19 ? _GEN_293 : _GEN_193; // @[IssueArbiter.scala 107:70]
  wire  _GEN_344 = issue_valid_0 & _T_19 ? _GEN_294 : _GEN_194; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_345 = issue_valid_0 & _T_19 ? _GEN_295 : _GEN_195; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_346 = issue_valid_0 & _T_19 ? _GEN_296 : _GEN_196; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_351 = issue_valid_0 & _T_19 ? _GEN_301 : _GEN_201; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_352 = issue_valid_0 & _T_19 ? _GEN_302 : _GEN_202; // @[IssueArbiter.scala 107:70]
  wire  _GEN_354 = issue_valid_0 & _T_19 ? _GEN_304 : _GEN_204; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_355 = ~mdu_occupy ? io_insts_in_1_inst : _GEN_330; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_356 = ~mdu_occupy ? io_insts_in_1_ysyx_print : _GEN_331; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [31:0] _GEN_360 = ~mdu_occupy ? io_insts_in_1_pc : _GEN_335; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [19:0] _GEN_361 = ~mdu_occupy ? io_insts_in_1_imm : _GEN_336; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_362 = ~mdu_occupy ? io_insts_in_1_rd : _GEN_337; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_367 = ~mdu_occupy ? io_insts_in_1_alu_expand : _GEN_342; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_368 = ~mdu_occupy ? io_insts_in_1_alu_op : _GEN_343; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_369 = ~mdu_occupy ? io_insts_in_1_write_dest : _GEN_344; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_370 = ~mdu_occupy ? io_insts_in_1_src_b : _GEN_345; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_371 = ~mdu_occupy ? io_insts_in_1_src_a : _GEN_346; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [63:0] _GEN_376 = ~mdu_occupy ? io_rss_in_1 : _GEN_351; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 116:25]
  wire [63:0] _GEN_377 = ~mdu_occupy ? io_rts_in_1 : _GEN_352; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 117:25]
  wire  _GEN_379 = ~mdu_occupy | _GEN_354; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 119:32]
  wire [31:0] _GEN_380 = ~alu_occupy ? io_insts_in_1_inst : _GEN_305; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_381 = ~alu_occupy ? io_insts_in_1_ysyx_print : _GEN_306; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_382 = ~alu_occupy ? io_insts_in_1_ysyx_debug : _GEN_307; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_383 = ~alu_occupy ? io_insts_in_1_target_pc : _GEN_308; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_384 = ~alu_occupy ? io_insts_in_1_predict_taken : _GEN_309; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_385 = ~alu_occupy ? io_insts_in_1_pc : _GEN_310; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [19:0] _GEN_386 = ~alu_occupy ? io_insts_in_1_imm : _GEN_311; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_387 = ~alu_occupy ? io_insts_in_1_rd : _GEN_312; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_389 = ~alu_occupy ? io_insts_in_1_rs1 : _GEN_314; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_390 = ~alu_occupy ? io_insts_in_1_write_src : _GEN_315; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_392 = ~alu_occupy ? io_insts_in_1_alu_expand : _GEN_317; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_393 = ~alu_occupy ? io_insts_in_1_alu_op : _GEN_318; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_394 = ~alu_occupy ? io_insts_in_1_write_dest : _GEN_319; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_395 = ~alu_occupy ? io_insts_in_1_src_b : _GEN_320; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_396 = ~alu_occupy ? io_insts_in_1_src_a : _GEN_321; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_397 = ~alu_occupy ? io_insts_in_1_branch_type : _GEN_322; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_398 = ~alu_occupy ? io_insts_in_1_alu_mdu_lsu : _GEN_323; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_399 = ~alu_occupy ? io_insts_in_1_next_pc : _GEN_324; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_400 = ~alu_occupy ? io_insts_in_1_illegal : _GEN_325; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [63:0] _GEN_401 = ~alu_occupy ? io_rss_in_1 : _GEN_326; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 110:25]
  wire [63:0] _GEN_402 = ~alu_occupy ? io_rts_in_1 : _GEN_327; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 111:25]
  wire  _GEN_404 = ~alu_occupy | _GEN_329; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 113:32]
  wire [31:0] _GEN_405 = ~alu_occupy ? _GEN_330 : _GEN_355; // @[IssueArbiter.scala 108:27]
  wire  _GEN_406 = ~alu_occupy ? _GEN_331 : _GEN_356; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_410 = ~alu_occupy ? _GEN_335 : _GEN_360; // @[IssueArbiter.scala 108:27]
  wire [19:0] _GEN_411 = ~alu_occupy ? _GEN_336 : _GEN_361; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_412 = ~alu_occupy ? _GEN_337 : _GEN_362; // @[IssueArbiter.scala 108:27]
  wire  _GEN_417 = ~alu_occupy ? _GEN_342 : _GEN_367; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_418 = ~alu_occupy ? _GEN_343 : _GEN_368; // @[IssueArbiter.scala 108:27]
  wire  _GEN_419 = ~alu_occupy ? _GEN_344 : _GEN_369; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_420 = ~alu_occupy ? _GEN_345 : _GEN_370; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_421 = ~alu_occupy ? _GEN_346 : _GEN_371; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_426 = ~alu_occupy ? _GEN_351 : _GEN_376; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_427 = ~alu_occupy ? _GEN_352 : _GEN_377; // @[IssueArbiter.scala 108:27]
  wire  _GEN_428 = ~alu_occupy ? 1'h0 : _T_48; // @[IssueArbiter.scala 108:27]
  wire  _GEN_429 = ~alu_occupy ? _GEN_354 : _GEN_379; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_430 = issue_valid_1 & _T_20 ? _GEN_380 : _GEN_305; // @[IssueArbiter.scala 107:70]
  wire  _GEN_431 = issue_valid_1 & _T_20 ? _GEN_381 : _GEN_306; // @[IssueArbiter.scala 107:70]
  wire  _GEN_432 = issue_valid_1 & _T_20 ? _GEN_382 : _GEN_307; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_433 = issue_valid_1 & _T_20 ? _GEN_383 : _GEN_308; // @[IssueArbiter.scala 107:70]
  wire  _GEN_434 = issue_valid_1 & _T_20 ? _GEN_384 : _GEN_309; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_435 = issue_valid_1 & _T_20 ? _GEN_385 : _GEN_310; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_436 = issue_valid_1 & _T_20 ? _GEN_386 : _GEN_311; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_437 = issue_valid_1 & _T_20 ? _GEN_387 : _GEN_312; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_439 = issue_valid_1 & _T_20 ? _GEN_389 : _GEN_314; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_440 = issue_valid_1 & _T_20 ? _GEN_390 : _GEN_315; // @[IssueArbiter.scala 107:70]
  wire  _GEN_442 = issue_valid_1 & _T_20 ? _GEN_392 : _GEN_317; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_443 = issue_valid_1 & _T_20 ? _GEN_393 : _GEN_318; // @[IssueArbiter.scala 107:70]
  wire  _GEN_444 = issue_valid_1 & _T_20 ? _GEN_394 : _GEN_319; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_445 = issue_valid_1 & _T_20 ? _GEN_395 : _GEN_320; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_446 = issue_valid_1 & _T_20 ? _GEN_396 : _GEN_321; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_447 = issue_valid_1 & _T_20 ? _GEN_397 : _GEN_322; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_448 = issue_valid_1 & _T_20 ? _GEN_398 : _GEN_323; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_449 = issue_valid_1 & _T_20 ? _GEN_399 : _GEN_324; // @[IssueArbiter.scala 107:70]
  wire  _GEN_450 = issue_valid_1 & _T_20 ? _GEN_400 : _GEN_325; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_451 = issue_valid_1 & _T_20 ? _GEN_401 : _GEN_326; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_452 = issue_valid_1 & _T_20 ? _GEN_402 : _GEN_327; // @[IssueArbiter.scala 107:70]
  wire  _GEN_453 = issue_valid_1 & _T_20 & _T_47; // @[IssueArbiter.scala 107:70]
  wire  _GEN_454 = issue_valid_1 & _T_20 ? _GEN_404 : _GEN_329; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_455 = issue_valid_1 & _T_20 ? _GEN_405 : _GEN_330; // @[IssueArbiter.scala 107:70]
  wire  _GEN_456 = issue_valid_1 & _T_20 ? _GEN_406 : _GEN_331; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_460 = issue_valid_1 & _T_20 ? _GEN_410 : _GEN_335; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_461 = issue_valid_1 & _T_20 ? _GEN_411 : _GEN_336; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_462 = issue_valid_1 & _T_20 ? _GEN_412 : _GEN_337; // @[IssueArbiter.scala 107:70]
  wire  _GEN_467 = issue_valid_1 & _T_20 ? _GEN_417 : _GEN_342; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_468 = issue_valid_1 & _T_20 ? _GEN_418 : _GEN_343; // @[IssueArbiter.scala 107:70]
  wire  _GEN_469 = issue_valid_1 & _T_20 ? _GEN_419 : _GEN_344; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_470 = issue_valid_1 & _T_20 ? _GEN_420 : _GEN_345; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_471 = issue_valid_1 & _T_20 ? _GEN_421 : _GEN_346; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_476 = issue_valid_1 & _T_20 ? _GEN_426 : _GEN_351; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_477 = issue_valid_1 & _T_20 ? _GEN_427 : _GEN_352; // @[IssueArbiter.scala 107:70]
  wire  _GEN_478 = issue_valid_1 & _T_20 & _GEN_428; // @[IssueArbiter.scala 107:70]
  wire  _GEN_479 = issue_valid_1 & _T_20 ? _GEN_429 : _GEN_354; // @[IssueArbiter.scala 107:70]
  wire  _T_55 = 2'h2 == io_insts_in_1_alu_mdu_lsu; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_480 = _T_55 ? io_insts_in_1_inst : _GEN_205; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire  _GEN_481 = _T_55 ? io_insts_in_1_ysyx_print : _GEN_206; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [31:0] _GEN_485 = _T_55 ? io_insts_in_1_pc : _GEN_210; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [19:0] _GEN_486 = _T_55 ? io_insts_in_1_imm : _GEN_211; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [4:0] _GEN_487 = _T_55 ? io_insts_in_1_rd : _GEN_212; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [2:0] _GEN_491 = _T_55 ? io_insts_in_1_mem_width : _GEN_216; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [4:0] _GEN_493 = _T_55 ? io_insts_in_1_alu_op : _GEN_218; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire  _GEN_494 = _T_55 ? io_insts_in_1_write_dest : _GEN_219; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [1:0] _GEN_496 = _T_55 ? io_insts_in_1_src_a : _GEN_221; // @[Conditional.scala 39:67 IssueArbiter.scala 97:27]
  wire [63:0] _GEN_501 = _T_55 ? io_rss_in_1 : _GEN_226; // @[Conditional.scala 39:67 IssueArbiter.scala 98:25]
  wire [63:0] _GEN_502 = _T_55 ? io_rts_in_1 : _GEN_227; // @[Conditional.scala 39:67 IssueArbiter.scala 99:25]
  wire  _GEN_504 = _T_55 | _GEN_229; // @[Conditional.scala 39:67 IssueArbiter.scala 101:32]
  wire [31:0] _GEN_505 = _T_54 ? io_insts_in_1_inst : _GEN_455; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire  _GEN_506 = _T_54 ? io_insts_in_1_ysyx_print : _GEN_456; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [31:0] _GEN_510 = _T_54 ? io_insts_in_1_pc : _GEN_460; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [19:0] _GEN_511 = _T_54 ? io_insts_in_1_imm : _GEN_461; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [4:0] _GEN_512 = _T_54 ? io_insts_in_1_rd : _GEN_462; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire  _GEN_517 = _T_54 ? io_insts_in_1_alu_expand : _GEN_467; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [4:0] _GEN_518 = _T_54 ? io_insts_in_1_alu_op : _GEN_468; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire  _GEN_519 = _T_54 ? io_insts_in_1_write_dest : _GEN_469; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [1:0] _GEN_520 = _T_54 ? io_insts_in_1_src_b : _GEN_470; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [1:0] _GEN_521 = _T_54 ? io_insts_in_1_src_a : _GEN_471; // @[Conditional.scala 39:67 IssueArbiter.scala 89:27]
  wire [63:0] _GEN_526 = _T_54 ? io_rss_in_1 : _GEN_476; // @[Conditional.scala 39:67 IssueArbiter.scala 90:25]
  wire [63:0] _GEN_527 = _T_54 ? io_rts_in_1 : _GEN_477; // @[Conditional.scala 39:67 IssueArbiter.scala 91:25]
  wire  _GEN_528 = _T_54 | _GEN_478; // @[Conditional.scala 39:67 IssueArbiter.scala 92:29]
  wire  _GEN_529 = _T_54 | _GEN_479; // @[Conditional.scala 39:67 IssueArbiter.scala 93:32]
  wire [31:0] _GEN_531 = _T_54 ? _GEN_205 : _GEN_480; // @[Conditional.scala 39:67]
  wire  _GEN_532 = _T_54 ? _GEN_206 : _GEN_481; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_536 = _T_54 ? _GEN_210 : _GEN_485; // @[Conditional.scala 39:67]
  wire [19:0] _GEN_537 = _T_54 ? _GEN_211 : _GEN_486; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_538 = _T_54 ? _GEN_212 : _GEN_487; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_542 = _T_54 ? _GEN_216 : _GEN_491; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_544 = _T_54 ? _GEN_218 : _GEN_493; // @[Conditional.scala 39:67]
  wire  _GEN_545 = _T_54 ? _GEN_219 : _GEN_494; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_547 = _T_54 ? _GEN_221 : _GEN_496; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_552 = _T_54 ? _GEN_226 : _GEN_501; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_553 = _T_54 ? _GEN_227 : _GEN_502; // @[Conditional.scala 39:67]
  wire  _GEN_554 = _T_54 ? 1'h0 : _T_55; // @[Conditional.scala 39:67]
  wire  _GEN_555 = _T_54 ? _GEN_229 : _GEN_504; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_556 = _T_53 ? io_insts_in_1_inst : _GEN_430; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_557 = _T_53 ? io_insts_in_1_ysyx_print : _GEN_431; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_558 = _T_53 ? io_insts_in_1_ysyx_debug : _GEN_432; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [31:0] _GEN_559 = _T_53 ? io_insts_in_1_target_pc : _GEN_433; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_560 = _T_53 ? io_insts_in_1_predict_taken : _GEN_434; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [31:0] _GEN_561 = _T_53 ? io_insts_in_1_pc : _GEN_435; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [19:0] _GEN_562 = _T_53 ? io_insts_in_1_imm : _GEN_436; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [4:0] _GEN_563 = _T_53 ? io_insts_in_1_rd : _GEN_437; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [4:0] _GEN_565 = _T_53 ? io_insts_in_1_rs1 : _GEN_439; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [1:0] _GEN_566 = _T_53 ? io_insts_in_1_write_src : _GEN_440; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_568 = _T_53 ? io_insts_in_1_alu_expand : _GEN_442; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [4:0] _GEN_569 = _T_53 ? io_insts_in_1_alu_op : _GEN_443; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_570 = _T_53 ? io_insts_in_1_write_dest : _GEN_444; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [1:0] _GEN_571 = _T_53 ? io_insts_in_1_src_b : _GEN_445; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [1:0] _GEN_572 = _T_53 ? io_insts_in_1_src_a : _GEN_446; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [3:0] _GEN_573 = _T_53 ? io_insts_in_1_branch_type : _GEN_447; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [1:0] _GEN_574 = _T_53 ? io_insts_in_1_alu_mdu_lsu : _GEN_448; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [3:0] _GEN_575 = _T_53 ? io_insts_in_1_next_pc : _GEN_449; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire  _GEN_576 = _T_53 ? io_insts_in_1_illegal : _GEN_450; // @[Conditional.scala 40:58 IssueArbiter.scala 81:27]
  wire [63:0] _GEN_577 = _T_53 ? io_rss_in_1 : _GEN_451; // @[Conditional.scala 40:58 IssueArbiter.scala 82:25]
  wire [63:0] _GEN_578 = _T_53 ? io_rts_in_1 : _GEN_452; // @[Conditional.scala 40:58 IssueArbiter.scala 83:25]
  wire  _GEN_579 = _T_53 | _GEN_453; // @[Conditional.scala 40:58 IssueArbiter.scala 84:29]
  wire  _GEN_580 = _T_53 | _GEN_454; // @[Conditional.scala 40:58 IssueArbiter.scala 85:32]
  wire [31:0] _GEN_582 = _T_53 ? _GEN_455 : _GEN_505; // @[Conditional.scala 40:58]
  wire  _GEN_583 = _T_53 ? _GEN_456 : _GEN_506; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_587 = _T_53 ? _GEN_460 : _GEN_510; // @[Conditional.scala 40:58]
  wire [19:0] _GEN_588 = _T_53 ? _GEN_461 : _GEN_511; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_589 = _T_53 ? _GEN_462 : _GEN_512; // @[Conditional.scala 40:58]
  wire  _GEN_594 = _T_53 ? _GEN_467 : _GEN_517; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_595 = _T_53 ? _GEN_468 : _GEN_518; // @[Conditional.scala 40:58]
  wire  _GEN_596 = _T_53 ? _GEN_469 : _GEN_519; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_597 = _T_53 ? _GEN_470 : _GEN_520; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_598 = _T_53 ? _GEN_471 : _GEN_521; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_603 = _T_53 ? _GEN_476 : _GEN_526; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_604 = _T_53 ? _GEN_477 : _GEN_527; // @[Conditional.scala 40:58]
  wire  _GEN_605 = _T_53 ? _GEN_478 : _GEN_528; // @[Conditional.scala 40:58]
  wire  _GEN_606 = _T_53 ? _GEN_479 : _GEN_529; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_608 = _T_53 ? _GEN_205 : _GEN_531; // @[Conditional.scala 40:58]
  wire  _GEN_609 = _T_53 ? _GEN_206 : _GEN_532; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_613 = _T_53 ? _GEN_210 : _GEN_536; // @[Conditional.scala 40:58]
  wire [19:0] _GEN_614 = _T_53 ? _GEN_211 : _GEN_537; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_615 = _T_53 ? _GEN_212 : _GEN_538; // @[Conditional.scala 40:58]
  wire [2:0] _GEN_619 = _T_53 ? _GEN_216 : _GEN_542; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_621 = _T_53 ? _GEN_218 : _GEN_544; // @[Conditional.scala 40:58]
  wire  _GEN_622 = _T_53 ? _GEN_219 : _GEN_545; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_624 = _T_53 ? _GEN_221 : _GEN_547; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_629 = _T_53 ? _GEN_226 : _GEN_552; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_630 = _T_53 ? _GEN_227 : _GEN_553; // @[Conditional.scala 40:58]
  wire  _GEN_631 = _T_53 ? 1'h0 : _GEN_554; // @[Conditional.scala 40:58]
  wire  _GEN_632 = _T_53 ? _GEN_229 : _GEN_555; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_633 = issue_valid_1 ? _GEN_556 : _GEN_430; // @[IssueArbiter.scala 78:26]
  wire  _GEN_634 = issue_valid_1 ? _GEN_557 : _GEN_431; // @[IssueArbiter.scala 78:26]
  wire  _GEN_635 = issue_valid_1 ? _GEN_558 : _GEN_432; // @[IssueArbiter.scala 78:26]
  wire [31:0] _GEN_636 = issue_valid_1 ? _GEN_559 : _GEN_433; // @[IssueArbiter.scala 78:26]
  wire  _GEN_637 = issue_valid_1 ? _GEN_560 : _GEN_434; // @[IssueArbiter.scala 78:26]
  wire [31:0] _GEN_638 = issue_valid_1 ? _GEN_561 : _GEN_435; // @[IssueArbiter.scala 78:26]
  wire [19:0] _GEN_639 = issue_valid_1 ? _GEN_562 : _GEN_436; // @[IssueArbiter.scala 78:26]
  wire [4:0] _GEN_640 = issue_valid_1 ? _GEN_563 : _GEN_437; // @[IssueArbiter.scala 78:26]
  wire [4:0] _GEN_642 = issue_valid_1 ? _GEN_565 : _GEN_439; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_643 = issue_valid_1 ? _GEN_566 : _GEN_440; // @[IssueArbiter.scala 78:26]
  wire  _GEN_645 = issue_valid_1 ? _GEN_568 : _GEN_442; // @[IssueArbiter.scala 78:26]
  wire [4:0] _GEN_646 = issue_valid_1 ? _GEN_569 : _GEN_443; // @[IssueArbiter.scala 78:26]
  wire  _GEN_647 = issue_valid_1 ? _GEN_570 : _GEN_444; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_648 = issue_valid_1 ? _GEN_571 : _GEN_445; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_649 = issue_valid_1 ? _GEN_572 : _GEN_446; // @[IssueArbiter.scala 78:26]
  wire [3:0] _GEN_650 = issue_valid_1 ? _GEN_573 : _GEN_447; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_651 = issue_valid_1 ? _GEN_574 : _GEN_448; // @[IssueArbiter.scala 78:26]
  wire [3:0] _GEN_652 = issue_valid_1 ? _GEN_575 : _GEN_449; // @[IssueArbiter.scala 78:26]
  wire  _GEN_653 = issue_valid_1 ? _GEN_576 : _GEN_450; // @[IssueArbiter.scala 78:26]
  wire [63:0] _GEN_654 = issue_valid_1 ? _GEN_577 : _GEN_451; // @[IssueArbiter.scala 78:26]
  wire [63:0] _GEN_655 = issue_valid_1 ? _GEN_578 : _GEN_452; // @[IssueArbiter.scala 78:26]
  wire  _GEN_656 = issue_valid_1 ? _GEN_579 : _GEN_453; // @[IssueArbiter.scala 78:26]
  wire  _GEN_657 = issue_valid_1 ? _GEN_580 : _GEN_454; // @[IssueArbiter.scala 78:26]
  wire [31:0] _GEN_659 = issue_valid_1 ? _GEN_582 : _GEN_455; // @[IssueArbiter.scala 78:26]
  wire  _GEN_660 = issue_valid_1 ? _GEN_583 : _GEN_456; // @[IssueArbiter.scala 78:26]
  wire [31:0] _GEN_664 = issue_valid_1 ? _GEN_587 : _GEN_460; // @[IssueArbiter.scala 78:26]
  wire [19:0] _GEN_665 = issue_valid_1 ? _GEN_588 : _GEN_461; // @[IssueArbiter.scala 78:26]
  wire [4:0] _GEN_666 = issue_valid_1 ? _GEN_589 : _GEN_462; // @[IssueArbiter.scala 78:26]
  wire  _GEN_671 = issue_valid_1 ? _GEN_594 : _GEN_467; // @[IssueArbiter.scala 78:26]
  wire [4:0] _GEN_672 = issue_valid_1 ? _GEN_595 : _GEN_468; // @[IssueArbiter.scala 78:26]
  wire  _GEN_673 = issue_valid_1 ? _GEN_596 : _GEN_469; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_674 = issue_valid_1 ? _GEN_597 : _GEN_470; // @[IssueArbiter.scala 78:26]
  wire [1:0] _GEN_675 = issue_valid_1 ? _GEN_598 : _GEN_471; // @[IssueArbiter.scala 78:26]
  wire [63:0] _GEN_680 = issue_valid_1 ? _GEN_603 : _GEN_476; // @[IssueArbiter.scala 78:26]
  wire [63:0] _GEN_681 = issue_valid_1 ? _GEN_604 : _GEN_477; // @[IssueArbiter.scala 78:26]
  wire  _GEN_682 = issue_valid_1 ? _GEN_605 : _GEN_478; // @[IssueArbiter.scala 78:26]
  wire  _GEN_683 = issue_valid_1 ? _GEN_606 : _GEN_479; // @[IssueArbiter.scala 78:26]
  wire  _GEN_708 = issue_valid_1 & _GEN_631; // @[IssueArbiter.scala 78:26]
  wire [31:0] _GEN_710 = ~mdu_occupy ? io_insts_in_0_inst : _GEN_659; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_711 = ~mdu_occupy ? io_insts_in_0_ysyx_print : _GEN_660; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [31:0] _GEN_715 = ~mdu_occupy ? io_insts_in_0_pc : _GEN_664; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [19:0] _GEN_716 = ~mdu_occupy ? io_insts_in_0_imm : _GEN_665; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_717 = ~mdu_occupy ? io_insts_in_0_rd : _GEN_666; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_722 = ~mdu_occupy ? io_insts_in_0_alu_expand : _GEN_671; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_723 = ~mdu_occupy ? io_insts_in_0_alu_op : _GEN_672; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_724 = ~mdu_occupy ? io_insts_in_0_write_dest : _GEN_673; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_725 = ~mdu_occupy ? io_insts_in_0_src_b : _GEN_674; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_726 = ~mdu_occupy ? io_insts_in_0_src_a : _GEN_675; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [63:0] _GEN_731 = ~mdu_occupy ? io_rss_in_0 : _GEN_680; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 116:25]
  wire [63:0] _GEN_732 = ~mdu_occupy ? io_rts_in_0 : _GEN_681; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 117:25]
  wire  _GEN_733 = ~mdu_occupy ? 1'h0 : _GEN_682; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 118:29]
  wire  _GEN_734 = ~mdu_occupy | _GEN_683; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 119:32]
  wire [31:0] _GEN_735 = ~alu_occupy ? io_insts_in_0_inst : _GEN_633; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_736 = ~alu_occupy ? io_insts_in_0_ysyx_print : _GEN_634; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_737 = ~alu_occupy ? io_insts_in_0_ysyx_debug : _GEN_635; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_738 = ~alu_occupy ? io_insts_in_0_target_pc : _GEN_636; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_739 = ~alu_occupy ? io_insts_in_0_predict_taken : _GEN_637; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_740 = ~alu_occupy ? io_insts_in_0_pc : _GEN_638; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [19:0] _GEN_741 = ~alu_occupy ? io_insts_in_0_imm : _GEN_639; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_742 = ~alu_occupy ? io_insts_in_0_rd : _GEN_640; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_744 = ~alu_occupy ? io_insts_in_0_rs1 : _GEN_642; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_745 = ~alu_occupy ? io_insts_in_0_write_src : _GEN_643; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_747 = ~alu_occupy ? io_insts_in_0_alu_expand : _GEN_645; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_748 = ~alu_occupy ? io_insts_in_0_alu_op : _GEN_646; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_749 = ~alu_occupy ? io_insts_in_0_write_dest : _GEN_647; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_750 = ~alu_occupy ? io_insts_in_0_src_b : _GEN_648; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_751 = ~alu_occupy ? io_insts_in_0_src_a : _GEN_649; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_752 = ~alu_occupy ? io_insts_in_0_branch_type : _GEN_650; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_753 = ~alu_occupy ? io_insts_in_0_alu_mdu_lsu : _GEN_651; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_754 = ~alu_occupy ? io_insts_in_0_next_pc : _GEN_652; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_755 = ~alu_occupy ? io_insts_in_0_illegal : _GEN_653; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [63:0] _GEN_756 = ~alu_occupy ? io_rss_in_0 : _GEN_654; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 110:25]
  wire [63:0] _GEN_757 = ~alu_occupy ? io_rts_in_0 : _GEN_655; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 111:25]
  wire  _GEN_758 = ~alu_occupy ? 1'h0 : _GEN_656; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 112:29]
  wire  _GEN_759 = ~alu_occupy | _GEN_657; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 113:32]
  wire [31:0] _GEN_760 = ~alu_occupy ? _GEN_659 : _GEN_710; // @[IssueArbiter.scala 108:27]
  wire  _GEN_761 = ~alu_occupy ? _GEN_660 : _GEN_711; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_765 = ~alu_occupy ? _GEN_664 : _GEN_715; // @[IssueArbiter.scala 108:27]
  wire [19:0] _GEN_766 = ~alu_occupy ? _GEN_665 : _GEN_716; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_767 = ~alu_occupy ? _GEN_666 : _GEN_717; // @[IssueArbiter.scala 108:27]
  wire  _GEN_772 = ~alu_occupy ? _GEN_671 : _GEN_722; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_773 = ~alu_occupy ? _GEN_672 : _GEN_723; // @[IssueArbiter.scala 108:27]
  wire  _GEN_774 = ~alu_occupy ? _GEN_673 : _GEN_724; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_775 = ~alu_occupy ? _GEN_674 : _GEN_725; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_776 = ~alu_occupy ? _GEN_675 : _GEN_726; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_781 = ~alu_occupy ? _GEN_680 : _GEN_731; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_782 = ~alu_occupy ? _GEN_681 : _GEN_732; // @[IssueArbiter.scala 108:27]
  wire  _GEN_783 = ~alu_occupy ? _GEN_682 : _GEN_733; // @[IssueArbiter.scala 108:27]
  wire  _GEN_784 = ~alu_occupy ? _GEN_683 : _GEN_734; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_785 = issue_valid_0 & _T_19 ? _GEN_735 : _GEN_633; // @[IssueArbiter.scala 107:70]
  wire  _GEN_786 = issue_valid_0 & _T_19 ? _GEN_736 : _GEN_634; // @[IssueArbiter.scala 107:70]
  wire  _GEN_787 = issue_valid_0 & _T_19 ? _GEN_737 : _GEN_635; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_788 = issue_valid_0 & _T_19 ? _GEN_738 : _GEN_636; // @[IssueArbiter.scala 107:70]
  wire  _GEN_789 = issue_valid_0 & _T_19 ? _GEN_739 : _GEN_637; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_790 = issue_valid_0 & _T_19 ? _GEN_740 : _GEN_638; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_791 = issue_valid_0 & _T_19 ? _GEN_741 : _GEN_639; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_792 = issue_valid_0 & _T_19 ? _GEN_742 : _GEN_640; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_794 = issue_valid_0 & _T_19 ? _GEN_744 : _GEN_642; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_795 = issue_valid_0 & _T_19 ? _GEN_745 : _GEN_643; // @[IssueArbiter.scala 107:70]
  wire  _GEN_797 = issue_valid_0 & _T_19 ? _GEN_747 : _GEN_645; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_798 = issue_valid_0 & _T_19 ? _GEN_748 : _GEN_646; // @[IssueArbiter.scala 107:70]
  wire  _GEN_799 = issue_valid_0 & _T_19 ? _GEN_749 : _GEN_647; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_800 = issue_valid_0 & _T_19 ? _GEN_750 : _GEN_648; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_801 = issue_valid_0 & _T_19 ? _GEN_751 : _GEN_649; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_802 = issue_valid_0 & _T_19 ? _GEN_752 : _GEN_650; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_803 = issue_valid_0 & _T_19 ? _GEN_753 : _GEN_651; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_804 = issue_valid_0 & _T_19 ? _GEN_754 : _GEN_652; // @[IssueArbiter.scala 107:70]
  wire  _GEN_805 = issue_valid_0 & _T_19 ? _GEN_755 : _GEN_653; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_806 = issue_valid_0 & _T_19 ? _GEN_756 : _GEN_654; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_807 = issue_valid_0 & _T_19 ? _GEN_757 : _GEN_655; // @[IssueArbiter.scala 107:70]
  wire  _GEN_808 = issue_valid_0 & _T_19 ? _GEN_758 : _GEN_656; // @[IssueArbiter.scala 107:70]
  wire  _GEN_809 = issue_valid_0 & _T_19 ? _GEN_759 : _GEN_657; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_810 = issue_valid_0 & _T_19 ? _GEN_760 : _GEN_659; // @[IssueArbiter.scala 107:70]
  wire  _GEN_811 = issue_valid_0 & _T_19 ? _GEN_761 : _GEN_660; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_815 = issue_valid_0 & _T_19 ? _GEN_765 : _GEN_664; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_816 = issue_valid_0 & _T_19 ? _GEN_766 : _GEN_665; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_817 = issue_valid_0 & _T_19 ? _GEN_767 : _GEN_666; // @[IssueArbiter.scala 107:70]
  wire  _GEN_822 = issue_valid_0 & _T_19 ? _GEN_772 : _GEN_671; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_823 = issue_valid_0 & _T_19 ? _GEN_773 : _GEN_672; // @[IssueArbiter.scala 107:70]
  wire  _GEN_824 = issue_valid_0 & _T_19 ? _GEN_774 : _GEN_673; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_825 = issue_valid_0 & _T_19 ? _GEN_775 : _GEN_674; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_826 = issue_valid_0 & _T_19 ? _GEN_776 : _GEN_675; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_831 = issue_valid_0 & _T_19 ? _GEN_781 : _GEN_680; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_832 = issue_valid_0 & _T_19 ? _GEN_782 : _GEN_681; // @[IssueArbiter.scala 107:70]
  wire  _GEN_833 = issue_valid_0 & _T_19 ? _GEN_783 : _GEN_682; // @[IssueArbiter.scala 107:70]
  wire  _GEN_834 = issue_valid_0 & _T_19 ? _GEN_784 : _GEN_683; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_835 = ~mdu_occupy ? io_insts_in_1_inst : _GEN_810; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_836 = ~mdu_occupy ? io_insts_in_1_ysyx_print : _GEN_811; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [31:0] _GEN_840 = ~mdu_occupy ? io_insts_in_1_pc : _GEN_815; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [19:0] _GEN_841 = ~mdu_occupy ? io_insts_in_1_imm : _GEN_816; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_842 = ~mdu_occupy ? io_insts_in_1_rd : _GEN_817; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_847 = ~mdu_occupy ? io_insts_in_1_alu_expand : _GEN_822; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [4:0] _GEN_848 = ~mdu_occupy ? io_insts_in_1_alu_op : _GEN_823; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire  _GEN_849 = ~mdu_occupy ? io_insts_in_1_write_dest : _GEN_824; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_850 = ~mdu_occupy ? io_insts_in_1_src_b : _GEN_825; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [1:0] _GEN_851 = ~mdu_occupy ? io_insts_in_1_src_a : _GEN_826; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 115:27]
  wire [63:0] _GEN_856 = ~mdu_occupy ? io_rss_in_1 : _GEN_831; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 116:25]
  wire [63:0] _GEN_857 = ~mdu_occupy ? io_rts_in_1 : _GEN_832; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 117:25]
  wire  _GEN_858 = ~mdu_occupy | _GEN_833; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 118:29]
  wire  _GEN_859 = ~mdu_occupy | _GEN_834; // @[IssueArbiter.scala 114:34 IssueArbiter.scala 119:32]
  wire [31:0] _GEN_860 = ~alu_occupy ? io_insts_in_1_inst : _GEN_785; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_861 = ~alu_occupy ? io_insts_in_1_ysyx_print : _GEN_786; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_862 = ~alu_occupy ? io_insts_in_1_ysyx_debug : _GEN_787; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_863 = ~alu_occupy ? io_insts_in_1_target_pc : _GEN_788; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_864 = ~alu_occupy ? io_insts_in_1_predict_taken : _GEN_789; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [31:0] _GEN_865 = ~alu_occupy ? io_insts_in_1_pc : _GEN_790; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [19:0] _GEN_866 = ~alu_occupy ? io_insts_in_1_imm : _GEN_791; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_867 = ~alu_occupy ? io_insts_in_1_rd : _GEN_792; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_869 = ~alu_occupy ? io_insts_in_1_rs1 : _GEN_794; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_870 = ~alu_occupy ? io_insts_in_1_write_src : _GEN_795; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_872 = ~alu_occupy ? io_insts_in_1_alu_expand : _GEN_797; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [4:0] _GEN_873 = ~alu_occupy ? io_insts_in_1_alu_op : _GEN_798; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_874 = ~alu_occupy ? io_insts_in_1_write_dest : _GEN_799; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_875 = ~alu_occupy ? io_insts_in_1_src_b : _GEN_800; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_876 = ~alu_occupy ? io_insts_in_1_src_a : _GEN_801; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_877 = ~alu_occupy ? io_insts_in_1_branch_type : _GEN_802; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [1:0] _GEN_878 = ~alu_occupy ? io_insts_in_1_alu_mdu_lsu : _GEN_803; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [3:0] _GEN_879 = ~alu_occupy ? io_insts_in_1_next_pc : _GEN_804; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire  _GEN_880 = ~alu_occupy ? io_insts_in_1_illegal : _GEN_805; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 109:27]
  wire [63:0] _GEN_881 = ~alu_occupy ? io_rss_in_1 : _GEN_806; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 110:25]
  wire [63:0] _GEN_882 = ~alu_occupy ? io_rts_in_1 : _GEN_807; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 111:25]
  wire  _GEN_883 = ~alu_occupy | _GEN_808; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 112:29]
  wire  _GEN_884 = ~alu_occupy | _GEN_809; // @[IssueArbiter.scala 108:27 IssueArbiter.scala 113:32]
  wire [31:0] _GEN_885 = ~alu_occupy ? _GEN_810 : _GEN_835; // @[IssueArbiter.scala 108:27]
  wire  _GEN_886 = ~alu_occupy ? _GEN_811 : _GEN_836; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_890 = ~alu_occupy ? _GEN_815 : _GEN_840; // @[IssueArbiter.scala 108:27]
  wire [19:0] _GEN_891 = ~alu_occupy ? _GEN_816 : _GEN_841; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_892 = ~alu_occupy ? _GEN_817 : _GEN_842; // @[IssueArbiter.scala 108:27]
  wire  _GEN_897 = ~alu_occupy ? _GEN_822 : _GEN_847; // @[IssueArbiter.scala 108:27]
  wire [4:0] _GEN_898 = ~alu_occupy ? _GEN_823 : _GEN_848; // @[IssueArbiter.scala 108:27]
  wire  _GEN_899 = ~alu_occupy ? _GEN_824 : _GEN_849; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_900 = ~alu_occupy ? _GEN_825 : _GEN_850; // @[IssueArbiter.scala 108:27]
  wire [1:0] _GEN_901 = ~alu_occupy ? _GEN_826 : _GEN_851; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_906 = ~alu_occupy ? _GEN_831 : _GEN_856; // @[IssueArbiter.scala 108:27]
  wire [63:0] _GEN_907 = ~alu_occupy ? _GEN_832 : _GEN_857; // @[IssueArbiter.scala 108:27]
  wire  _GEN_908 = ~alu_occupy ? _GEN_833 : _GEN_858; // @[IssueArbiter.scala 108:27]
  wire  _GEN_909 = ~alu_occupy ? _GEN_834 : _GEN_859; // @[IssueArbiter.scala 108:27]
  wire [31:0] _GEN_910 = issue_valid_1 & _T_20 ? _GEN_860 : _GEN_785; // @[IssueArbiter.scala 107:70]
  wire  _GEN_911 = issue_valid_1 & _T_20 ? _GEN_861 : _GEN_786; // @[IssueArbiter.scala 107:70]
  wire  _GEN_912 = issue_valid_1 & _T_20 ? _GEN_862 : _GEN_787; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_913 = issue_valid_1 & _T_20 ? _GEN_863 : _GEN_788; // @[IssueArbiter.scala 107:70]
  wire  _GEN_914 = issue_valid_1 & _T_20 ? _GEN_864 : _GEN_789; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_915 = issue_valid_1 & _T_20 ? _GEN_865 : _GEN_790; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_916 = issue_valid_1 & _T_20 ? _GEN_866 : _GEN_791; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_917 = issue_valid_1 & _T_20 ? _GEN_867 : _GEN_792; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_919 = issue_valid_1 & _T_20 ? _GEN_869 : _GEN_794; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_920 = issue_valid_1 & _T_20 ? _GEN_870 : _GEN_795; // @[IssueArbiter.scala 107:70]
  wire  _GEN_922 = issue_valid_1 & _T_20 ? _GEN_872 : _GEN_797; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_923 = issue_valid_1 & _T_20 ? _GEN_873 : _GEN_798; // @[IssueArbiter.scala 107:70]
  wire  _GEN_924 = issue_valid_1 & _T_20 ? _GEN_874 : _GEN_799; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_925 = issue_valid_1 & _T_20 ? _GEN_875 : _GEN_800; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_926 = issue_valid_1 & _T_20 ? _GEN_876 : _GEN_801; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_927 = issue_valid_1 & _T_20 ? _GEN_877 : _GEN_802; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_928 = issue_valid_1 & _T_20 ? _GEN_878 : _GEN_803; // @[IssueArbiter.scala 107:70]
  wire [3:0] _GEN_929 = issue_valid_1 & _T_20 ? _GEN_879 : _GEN_804; // @[IssueArbiter.scala 107:70]
  wire  _GEN_930 = issue_valid_1 & _T_20 ? _GEN_880 : _GEN_805; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_931 = issue_valid_1 & _T_20 ? _GEN_881 : _GEN_806; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_932 = issue_valid_1 & _T_20 ? _GEN_882 : _GEN_807; // @[IssueArbiter.scala 107:70]
  wire  _GEN_933 = issue_valid_1 & _T_20 ? _GEN_883 : _GEN_808; // @[IssueArbiter.scala 107:70]
  wire  _GEN_934 = issue_valid_1 & _T_20 ? _GEN_884 : _GEN_809; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_935 = issue_valid_1 & _T_20 ? _GEN_885 : _GEN_810; // @[IssueArbiter.scala 107:70]
  wire  _GEN_936 = issue_valid_1 & _T_20 ? _GEN_886 : _GEN_811; // @[IssueArbiter.scala 107:70]
  wire [31:0] _GEN_940 = issue_valid_1 & _T_20 ? _GEN_890 : _GEN_815; // @[IssueArbiter.scala 107:70]
  wire [19:0] _GEN_941 = issue_valid_1 & _T_20 ? _GEN_891 : _GEN_816; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_942 = issue_valid_1 & _T_20 ? _GEN_892 : _GEN_817; // @[IssueArbiter.scala 107:70]
  wire  _GEN_947 = issue_valid_1 & _T_20 ? _GEN_897 : _GEN_822; // @[IssueArbiter.scala 107:70]
  wire [4:0] _GEN_948 = issue_valid_1 & _T_20 ? _GEN_898 : _GEN_823; // @[IssueArbiter.scala 107:70]
  wire  _GEN_949 = issue_valid_1 & _T_20 ? _GEN_899 : _GEN_824; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_950 = issue_valid_1 & _T_20 ? _GEN_900 : _GEN_825; // @[IssueArbiter.scala 107:70]
  wire [1:0] _GEN_951 = issue_valid_1 & _T_20 ? _GEN_901 : _GEN_826; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_956 = issue_valid_1 & _T_20 ? _GEN_906 : _GEN_831; // @[IssueArbiter.scala 107:70]
  wire [63:0] _GEN_957 = issue_valid_1 & _T_20 ? _GEN_907 : _GEN_832; // @[IssueArbiter.scala 107:70]
  wire  _GEN_958 = issue_valid_1 & _T_20 ? _GEN_908 : _GEN_833; // @[IssueArbiter.scala 107:70]
  wire  _GEN_959 = issue_valid_1 & _T_20 ? _GEN_909 : _GEN_834; // @[IssueArbiter.scala 107:70]
  wire  _GEN_983 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ? 1'h0 :
    _GEN_933; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 166:25]
  wire  _GEN_1008 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu | _GEN_958; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 171:25]
  assign io_rss_out_0 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_rss_in_0 : _GEN_931; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 164:21]
  assign io_rss_out_1 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_rss_in_1 : _GEN_956; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 169:21]
  assign io_rss_out_2 = issue_valid_1 ? _GEN_629 : _GEN_226; // @[IssueArbiter.scala 78:26]
  assign io_rts_out_0 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_rts_in_0 : _GEN_932; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 165:21]
  assign io_rts_out_1 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_rts_in_1 : _GEN_957; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 170:21]
  assign io_rts_out_2 = issue_valid_1 ? _GEN_630 : _GEN_227; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_0_illegal = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_0_illegal : _GEN_930; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_next_pc = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_0_next_pc : _GEN_929; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_alu_mdu_lsu = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_alu_mdu_lsu : _GEN_928; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_branch_type = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_branch_type : _GEN_927; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_src_a = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_0_src_a : _GEN_926; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_src_b = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_0_src_b : _GEN_925; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_write_dest = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_write_dest : _GEN_924; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_alu_op = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_0_alu_op : _GEN_923; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_alu_expand = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_alu_expand : _GEN_922; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_write_src = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_write_src : _GEN_920; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_rs1 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_0_rs1 : _GEN_919; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_rd = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_0_rd : _GEN_917; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_imm = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_0_imm : _GEN_916; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_pc = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_0_pc : _GEN_915; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_predict_taken = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_predict_taken : _GEN_914; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_target_pc = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_target_pc : _GEN_913; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_ysyx_debug = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_ysyx_debug : _GEN_912; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_ysyx_print = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_0_ysyx_print : _GEN_911; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_0_inst = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_0_inst : _GEN_910; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 163:23]
  assign io_insts_out_1_src_a = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_1_src_a : _GEN_951; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_src_b = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_1_src_b : _GEN_950; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_write_dest = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_1_write_dest : _GEN_949; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_alu_op = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu
     ? io_insts_in_1_alu_op : _GEN_948; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_alu_expand = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_1_alu_expand : _GEN_947; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_rd = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_1_rd : _GEN_942; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_imm = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_1_imm : _GEN_941; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_pc = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_1_pc : _GEN_940; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_ysyx_print = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu ==
    io_insts_in_1_alu_mdu_lsu ? io_insts_in_1_ysyx_print : _GEN_936; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_1_inst = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu ?
    io_insts_in_1_inst : _GEN_935; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 168:23]
  assign io_insts_out_2_src_a = issue_valid_1 ? _GEN_624 : _GEN_221; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_write_dest = issue_valid_1 ? _GEN_622 : _GEN_219; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_alu_op = issue_valid_1 ? _GEN_621 : _GEN_218; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_mem_width = issue_valid_1 ? _GEN_619 : _GEN_216; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_rd = issue_valid_1 ? _GEN_615 : _GEN_212; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_imm = issue_valid_1 ? _GEN_614 : _GEN_211; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_pc = issue_valid_1 ? _GEN_613 : _GEN_210; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_ysyx_print = issue_valid_1 ? _GEN_609 : _GEN_206; // @[IssueArbiter.scala 78:26]
  assign io_insts_out_2_inst = issue_valid_1 ? _GEN_608 : _GEN_205; // @[IssueArbiter.scala 78:26]
  assign io_issue_num = issue_valid_0 ? _GEN_1 : 2'h0; // @[IssueArbiter.scala 53:83 IssueArbiter.scala 52:16]
  assign io_issue_fu_valid_0 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu |
    _GEN_934; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 167:28]
  assign io_issue_fu_valid_1 = issue_valid_0 & issue_valid_1 & io_insts_in_0_alu_mdu_lsu == io_insts_in_1_alu_mdu_lsu |
    _GEN_959; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 172:28]
  assign io_issue_fu_valid_2 = issue_valid_1 ? _GEN_632 : _GEN_229; // @[IssueArbiter.scala 78:26]
  assign io_insts_order_0 = {{1'd0}, _GEN_983}; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 166:25]
  assign io_insts_order_1 = {{1'd0}, _GEN_1008}; // @[IssueArbiter.scala 162:105 IssueArbiter.scala 171:25]
  assign io_insts_order_2 = {{1'd0}, _GEN_708}; // @[IssueArbiter.scala 78:26]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs_addr_vec_0,
  input  [4:0]  io_rs_addr_vec_1,
  input  [4:0]  io_rs_addr_vec_2,
  input  [4:0]  io_rs_addr_vec_3,
  output [63:0] io_rs_data_vec_0,
  output [63:0] io_rs_data_vec_1,
  output [63:0] io_rs_data_vec_2,
  output [63:0] io_rs_data_vec_3,
  input         io_wen_vec_0,
  input         io_wen_vec_1,
  input  [4:0]  io_rd_addr_vec_0,
  input  [4:0]  io_rd_addr_vec_1,
  input  [63:0] io_rd_data_vec_0,
  input  [63:0] io_rd_data_vec_1,
  input  [4:0]  difftestSaddr,
  output [63:0] _WIRE_0_0,
  output [63:0] _WIRE_0_1,
  output [63:0] _WIRE_0_2,
  output [63:0] _WIRE_0_3,
  output [63:0] _WIRE_0_4,
  output [63:0] _WIRE_0_5,
  output [63:0] _WIRE_0_6,
  output [63:0] _WIRE_0_7,
  output [63:0] _WIRE_0_8,
  output [63:0] _WIRE_0_9,
  output [63:0] _WIRE_0_10,
  output [63:0] _WIRE_0_11,
  output [63:0] _WIRE_0_12,
  output [63:0] _WIRE_0_13,
  output [63:0] _WIRE_0_14,
  output [63:0] _WIRE_0_15,
  output [63:0] _WIRE_0_16,
  output [63:0] _WIRE_0_17,
  output [63:0] _WIRE_0_18,
  output [63:0] _WIRE_0_19,
  output [63:0] _WIRE_0_20,
  output [63:0] _WIRE_0_21,
  output [63:0] _WIRE_0_22,
  output [63:0] _WIRE_0_23,
  output [63:0] _WIRE_0_24,
  output [63:0] _WIRE_0_25,
  output [63:0] _WIRE_0_26,
  output [63:0] _WIRE_0_27,
  output [63:0] _WIRE_0_28,
  output [63:0] _WIRE_0_29,
  output [63:0] _WIRE_0_30,
  output [63:0] _WIRE_0_31,
  input  [31:0] difftestSval,
  input         difftestSync
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[RegFile.scala 20:21]
  reg [63:0] regs_1; // @[RegFile.scala 20:21]
  reg [63:0] regs_2; // @[RegFile.scala 20:21]
  reg [63:0] regs_3; // @[RegFile.scala 20:21]
  reg [63:0] regs_4; // @[RegFile.scala 20:21]
  reg [63:0] regs_5; // @[RegFile.scala 20:21]
  reg [63:0] regs_6; // @[RegFile.scala 20:21]
  reg [63:0] regs_7; // @[RegFile.scala 20:21]
  reg [63:0] regs_8; // @[RegFile.scala 20:21]
  reg [63:0] regs_9; // @[RegFile.scala 20:21]
  reg [63:0] regs_10; // @[RegFile.scala 20:21]
  reg [63:0] regs_11; // @[RegFile.scala 20:21]
  reg [63:0] regs_12; // @[RegFile.scala 20:21]
  reg [63:0] regs_13; // @[RegFile.scala 20:21]
  reg [63:0] regs_14; // @[RegFile.scala 20:21]
  reg [63:0] regs_15; // @[RegFile.scala 20:21]
  reg [63:0] regs_16; // @[RegFile.scala 20:21]
  reg [63:0] regs_17; // @[RegFile.scala 20:21]
  reg [63:0] regs_18; // @[RegFile.scala 20:21]
  reg [63:0] regs_19; // @[RegFile.scala 20:21]
  reg [63:0] regs_20; // @[RegFile.scala 20:21]
  reg [63:0] regs_21; // @[RegFile.scala 20:21]
  reg [63:0] regs_22; // @[RegFile.scala 20:21]
  reg [63:0] regs_23; // @[RegFile.scala 20:21]
  reg [63:0] regs_24; // @[RegFile.scala 20:21]
  reg [63:0] regs_25; // @[RegFile.scala 20:21]
  reg [63:0] regs_26; // @[RegFile.scala 20:21]
  reg [63:0] regs_27; // @[RegFile.scala 20:21]
  reg [63:0] regs_28; // @[RegFile.scala 20:21]
  reg [63:0] regs_29; // @[RegFile.scala 20:21]
  reg [63:0] regs_30; // @[RegFile.scala 20:21]
  reg [63:0] regs_31; // @[RegFile.scala 20:21]
  wire [63:0] _GEN_0 = regs_0; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_1 = 5'h1 == io_rs_addr_vec_0 ? regs_1 : regs_0; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_2 = 5'h2 == io_rs_addr_vec_0 ? regs_2 : _GEN_1; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_3 = 5'h3 == io_rs_addr_vec_0 ? regs_3 : _GEN_2; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_4 = 5'h4 == io_rs_addr_vec_0 ? regs_4 : _GEN_3; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_5 = 5'h5 == io_rs_addr_vec_0 ? regs_5 : _GEN_4; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_6 = 5'h6 == io_rs_addr_vec_0 ? regs_6 : _GEN_5; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_7 = 5'h7 == io_rs_addr_vec_0 ? regs_7 : _GEN_6; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_8 = 5'h8 == io_rs_addr_vec_0 ? regs_8 : _GEN_7; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_9 = 5'h9 == io_rs_addr_vec_0 ? regs_9 : _GEN_8; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_10 = 5'ha == io_rs_addr_vec_0 ? regs_10 : _GEN_9; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_11 = 5'hb == io_rs_addr_vec_0 ? regs_11 : _GEN_10; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_12 = 5'hc == io_rs_addr_vec_0 ? regs_12 : _GEN_11; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_13 = 5'hd == io_rs_addr_vec_0 ? regs_13 : _GEN_12; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_14 = 5'he == io_rs_addr_vec_0 ? regs_14 : _GEN_13; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_15 = 5'hf == io_rs_addr_vec_0 ? regs_15 : _GEN_14; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_16 = 5'h10 == io_rs_addr_vec_0 ? regs_16 : _GEN_15; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_17 = 5'h11 == io_rs_addr_vec_0 ? regs_17 : _GEN_16; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_18 = 5'h12 == io_rs_addr_vec_0 ? regs_18 : _GEN_17; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_19 = 5'h13 == io_rs_addr_vec_0 ? regs_19 : _GEN_18; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_20 = 5'h14 == io_rs_addr_vec_0 ? regs_20 : _GEN_19; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_21 = 5'h15 == io_rs_addr_vec_0 ? regs_21 : _GEN_20; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_22 = 5'h16 == io_rs_addr_vec_0 ? regs_22 : _GEN_21; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_23 = 5'h17 == io_rs_addr_vec_0 ? regs_23 : _GEN_22; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_24 = 5'h18 == io_rs_addr_vec_0 ? regs_24 : _GEN_23; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_25 = 5'h19 == io_rs_addr_vec_0 ? regs_25 : _GEN_24; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_26 = 5'h1a == io_rs_addr_vec_0 ? regs_26 : _GEN_25; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_27 = 5'h1b == io_rs_addr_vec_0 ? regs_27 : _GEN_26; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_28 = 5'h1c == io_rs_addr_vec_0 ? regs_28 : _GEN_27; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_29 = 5'h1d == io_rs_addr_vec_0 ? regs_29 : _GEN_28; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_30 = 5'h1e == io_rs_addr_vec_0 ? regs_30 : _GEN_29; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_31 = 5'h1f == io_rs_addr_vec_0 ? regs_31 : _GEN_30; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_33 = 5'h1 == io_rs_addr_vec_1 ? regs_1 : regs_0; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_34 = 5'h2 == io_rs_addr_vec_1 ? regs_2 : _GEN_33; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_35 = 5'h3 == io_rs_addr_vec_1 ? regs_3 : _GEN_34; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_36 = 5'h4 == io_rs_addr_vec_1 ? regs_4 : _GEN_35; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_37 = 5'h5 == io_rs_addr_vec_1 ? regs_5 : _GEN_36; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_38 = 5'h6 == io_rs_addr_vec_1 ? regs_6 : _GEN_37; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_39 = 5'h7 == io_rs_addr_vec_1 ? regs_7 : _GEN_38; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_40 = 5'h8 == io_rs_addr_vec_1 ? regs_8 : _GEN_39; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_41 = 5'h9 == io_rs_addr_vec_1 ? regs_9 : _GEN_40; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_42 = 5'ha == io_rs_addr_vec_1 ? regs_10 : _GEN_41; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_43 = 5'hb == io_rs_addr_vec_1 ? regs_11 : _GEN_42; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_44 = 5'hc == io_rs_addr_vec_1 ? regs_12 : _GEN_43; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_45 = 5'hd == io_rs_addr_vec_1 ? regs_13 : _GEN_44; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_46 = 5'he == io_rs_addr_vec_1 ? regs_14 : _GEN_45; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_47 = 5'hf == io_rs_addr_vec_1 ? regs_15 : _GEN_46; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_48 = 5'h10 == io_rs_addr_vec_1 ? regs_16 : _GEN_47; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_49 = 5'h11 == io_rs_addr_vec_1 ? regs_17 : _GEN_48; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_50 = 5'h12 == io_rs_addr_vec_1 ? regs_18 : _GEN_49; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_51 = 5'h13 == io_rs_addr_vec_1 ? regs_19 : _GEN_50; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_52 = 5'h14 == io_rs_addr_vec_1 ? regs_20 : _GEN_51; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_53 = 5'h15 == io_rs_addr_vec_1 ? regs_21 : _GEN_52; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_54 = 5'h16 == io_rs_addr_vec_1 ? regs_22 : _GEN_53; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_55 = 5'h17 == io_rs_addr_vec_1 ? regs_23 : _GEN_54; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_56 = 5'h18 == io_rs_addr_vec_1 ? regs_24 : _GEN_55; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_57 = 5'h19 == io_rs_addr_vec_1 ? regs_25 : _GEN_56; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_58 = 5'h1a == io_rs_addr_vec_1 ? regs_26 : _GEN_57; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_59 = 5'h1b == io_rs_addr_vec_1 ? regs_27 : _GEN_58; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_60 = 5'h1c == io_rs_addr_vec_1 ? regs_28 : _GEN_59; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_61 = 5'h1d == io_rs_addr_vec_1 ? regs_29 : _GEN_60; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_62 = 5'h1e == io_rs_addr_vec_1 ? regs_30 : _GEN_61; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_63 = 5'h1f == io_rs_addr_vec_1 ? regs_31 : _GEN_62; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_65 = 5'h1 == io_rs_addr_vec_2 ? regs_1 : regs_0; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_66 = 5'h2 == io_rs_addr_vec_2 ? regs_2 : _GEN_65; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_67 = 5'h3 == io_rs_addr_vec_2 ? regs_3 : _GEN_66; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_68 = 5'h4 == io_rs_addr_vec_2 ? regs_4 : _GEN_67; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_69 = 5'h5 == io_rs_addr_vec_2 ? regs_5 : _GEN_68; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_70 = 5'h6 == io_rs_addr_vec_2 ? regs_6 : _GEN_69; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_71 = 5'h7 == io_rs_addr_vec_2 ? regs_7 : _GEN_70; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_72 = 5'h8 == io_rs_addr_vec_2 ? regs_8 : _GEN_71; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_73 = 5'h9 == io_rs_addr_vec_2 ? regs_9 : _GEN_72; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_74 = 5'ha == io_rs_addr_vec_2 ? regs_10 : _GEN_73; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_75 = 5'hb == io_rs_addr_vec_2 ? regs_11 : _GEN_74; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_76 = 5'hc == io_rs_addr_vec_2 ? regs_12 : _GEN_75; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_77 = 5'hd == io_rs_addr_vec_2 ? regs_13 : _GEN_76; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_78 = 5'he == io_rs_addr_vec_2 ? regs_14 : _GEN_77; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_79 = 5'hf == io_rs_addr_vec_2 ? regs_15 : _GEN_78; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_80 = 5'h10 == io_rs_addr_vec_2 ? regs_16 : _GEN_79; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_81 = 5'h11 == io_rs_addr_vec_2 ? regs_17 : _GEN_80; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_82 = 5'h12 == io_rs_addr_vec_2 ? regs_18 : _GEN_81; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_83 = 5'h13 == io_rs_addr_vec_2 ? regs_19 : _GEN_82; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_84 = 5'h14 == io_rs_addr_vec_2 ? regs_20 : _GEN_83; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_85 = 5'h15 == io_rs_addr_vec_2 ? regs_21 : _GEN_84; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_86 = 5'h16 == io_rs_addr_vec_2 ? regs_22 : _GEN_85; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_87 = 5'h17 == io_rs_addr_vec_2 ? regs_23 : _GEN_86; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_88 = 5'h18 == io_rs_addr_vec_2 ? regs_24 : _GEN_87; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_89 = 5'h19 == io_rs_addr_vec_2 ? regs_25 : _GEN_88; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_90 = 5'h1a == io_rs_addr_vec_2 ? regs_26 : _GEN_89; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_91 = 5'h1b == io_rs_addr_vec_2 ? regs_27 : _GEN_90; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_92 = 5'h1c == io_rs_addr_vec_2 ? regs_28 : _GEN_91; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_93 = 5'h1d == io_rs_addr_vec_2 ? regs_29 : _GEN_92; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_94 = 5'h1e == io_rs_addr_vec_2 ? regs_30 : _GEN_93; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_95 = 5'h1f == io_rs_addr_vec_2 ? regs_31 : _GEN_94; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_97 = 5'h1 == io_rs_addr_vec_3 ? regs_1 : regs_0; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_98 = 5'h2 == io_rs_addr_vec_3 ? regs_2 : _GEN_97; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_99 = 5'h3 == io_rs_addr_vec_3 ? regs_3 : _GEN_98; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_100 = 5'h4 == io_rs_addr_vec_3 ? regs_4 : _GEN_99; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_101 = 5'h5 == io_rs_addr_vec_3 ? regs_5 : _GEN_100; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_102 = 5'h6 == io_rs_addr_vec_3 ? regs_6 : _GEN_101; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_103 = 5'h7 == io_rs_addr_vec_3 ? regs_7 : _GEN_102; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_104 = 5'h8 == io_rs_addr_vec_3 ? regs_8 : _GEN_103; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_105 = 5'h9 == io_rs_addr_vec_3 ? regs_9 : _GEN_104; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_106 = 5'ha == io_rs_addr_vec_3 ? regs_10 : _GEN_105; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_107 = 5'hb == io_rs_addr_vec_3 ? regs_11 : _GEN_106; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_108 = 5'hc == io_rs_addr_vec_3 ? regs_12 : _GEN_107; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_109 = 5'hd == io_rs_addr_vec_3 ? regs_13 : _GEN_108; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_110 = 5'he == io_rs_addr_vec_3 ? regs_14 : _GEN_109; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_111 = 5'hf == io_rs_addr_vec_3 ? regs_15 : _GEN_110; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_112 = 5'h10 == io_rs_addr_vec_3 ? regs_16 : _GEN_111; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_113 = 5'h11 == io_rs_addr_vec_3 ? regs_17 : _GEN_112; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_114 = 5'h12 == io_rs_addr_vec_3 ? regs_18 : _GEN_113; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_115 = 5'h13 == io_rs_addr_vec_3 ? regs_19 : _GEN_114; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_116 = 5'h14 == io_rs_addr_vec_3 ? regs_20 : _GEN_115; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_117 = 5'h15 == io_rs_addr_vec_3 ? regs_21 : _GEN_116; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_118 = 5'h16 == io_rs_addr_vec_3 ? regs_22 : _GEN_117; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_119 = 5'h17 == io_rs_addr_vec_3 ? regs_23 : _GEN_118; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_120 = 5'h18 == io_rs_addr_vec_3 ? regs_24 : _GEN_119; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_121 = 5'h19 == io_rs_addr_vec_3 ? regs_25 : _GEN_120; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_122 = 5'h1a == io_rs_addr_vec_3 ? regs_26 : _GEN_121; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_123 = 5'h1b == io_rs_addr_vec_3 ? regs_27 : _GEN_122; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_124 = 5'h1c == io_rs_addr_vec_3 ? regs_28 : _GEN_123; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_125 = 5'h1d == io_rs_addr_vec_3 ? regs_29 : _GEN_124; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_126 = 5'h1e == io_rs_addr_vec_3 ? regs_30 : _GEN_125; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_127 = 5'h1f == io_rs_addr_vec_3 ? regs_31 : _GEN_126; // @[RegFile.scala 22:23 RegFile.scala 22:23]
  wire [63:0] _GEN_128 = 5'h0 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_0; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_129 = 5'h1 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_1; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_130 = 5'h2 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_2; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_131 = 5'h3 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_3; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_132 = 5'h4 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_4; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_133 = 5'h5 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_5; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_134 = 5'h6 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_6; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_135 = 5'h7 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_7; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_136 = 5'h8 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_8; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_137 = 5'h9 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_9; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_138 = 5'ha == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_10; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_139 = 5'hb == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_11; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_140 = 5'hc == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_12; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_141 = 5'hd == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_13; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_142 = 5'he == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_14; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_143 = 5'hf == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_15; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_144 = 5'h10 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_16; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_145 = 5'h11 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_17; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_146 = 5'h12 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_18; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_147 = 5'h13 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_19; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_148 = 5'h14 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_20; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_149 = 5'h15 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_21; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_150 = 5'h16 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_22; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_151 = 5'h17 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_23; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_152 = 5'h18 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_24; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_153 = 5'h19 == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_25; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_154 = 5'h1a == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_26; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_155 = 5'h1b == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_27; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_156 = 5'h1c == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_28; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_157 = 5'h1d == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_29; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_158 = 5'h1e == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_30; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_159 = 5'h1f == io_rd_addr_vec_0 ? io_rd_data_vec_0 : regs_31; // @[RegFile.scala 26:31 RegFile.scala 26:31 RegFile.scala 20:21]
  wire [63:0] _GEN_160 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_128 : regs_0; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_161 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_129 : regs_1; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_162 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_130 : regs_2; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_163 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_131 : regs_3; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_164 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_132 : regs_4; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_165 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_133 : regs_5; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_166 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_134 : regs_6; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_167 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_135 : regs_7; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_168 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_136 : regs_8; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_169 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_137 : regs_9; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_170 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_138 : regs_10; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_171 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_139 : regs_11; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_172 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_140 : regs_12; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_173 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_141 : regs_13; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_174 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_142 : regs_14; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_175 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_143 : regs_15; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_176 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_144 : regs_16; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_177 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_145 : regs_17; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_178 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_146 : regs_18; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_179 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_147 : regs_19; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_180 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_148 : regs_20; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_181 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_149 : regs_21; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_182 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_150 : regs_22; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_183 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_151 : regs_23; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_184 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_152 : regs_24; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_185 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_153 : regs_25; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_186 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_154 : regs_26; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_187 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_155 : regs_27; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_188 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_156 : regs_28; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_189 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_157 : regs_29; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_190 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_158 : regs_30; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_191 = io_wen_vec_0 & |io_rd_addr_vec_0 ? _GEN_159 : regs_31; // @[RegFile.scala 25:50 RegFile.scala 20:21]
  wire [63:0] _GEN_192 = 5'h0 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_160; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_193 = 5'h1 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_161; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_194 = 5'h2 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_162; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_195 = 5'h3 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_163; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_196 = 5'h4 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_164; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_197 = 5'h5 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_165; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_198 = 5'h6 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_166; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_199 = 5'h7 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_167; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_200 = 5'h8 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_168; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_201 = 5'h9 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_169; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_202 = 5'ha == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_170; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_203 = 5'hb == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_171; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_204 = 5'hc == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_172; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_205 = 5'hd == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_173; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_206 = 5'he == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_174; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_207 = 5'hf == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_175; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_208 = 5'h10 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_176; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_209 = 5'h11 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_177; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_210 = 5'h12 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_178; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_211 = 5'h13 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_179; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_212 = 5'h14 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_180; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_213 = 5'h15 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_181; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_214 = 5'h16 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_182; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_215 = 5'h17 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_183; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_216 = 5'h18 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_184; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_217 = 5'h19 == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_185; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_218 = 5'h1a == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_186; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_219 = 5'h1b == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_187; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_220 = 5'h1c == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_188; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_221 = 5'h1d == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_189; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_222 = 5'h1e == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_190; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_223 = 5'h1f == io_rd_addr_vec_1 ? io_rd_data_vec_1 : _GEN_191; // @[RegFile.scala 26:31 RegFile.scala 26:31]
  wire [63:0] _GEN_224 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_192 : _GEN_160; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_225 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_193 : _GEN_161; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_226 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_194 : _GEN_162; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_227 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_195 : _GEN_163; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_228 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_196 : _GEN_164; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_229 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_197 : _GEN_165; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_230 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_198 : _GEN_166; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_231 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_199 : _GEN_167; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_232 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_200 : _GEN_168; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_233 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_201 : _GEN_169; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_234 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_202 : _GEN_170; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_235 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_203 : _GEN_171; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_236 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_204 : _GEN_172; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_237 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_205 : _GEN_173; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_238 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_206 : _GEN_174; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_239 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_207 : _GEN_175; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_240 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_208 : _GEN_176; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_241 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_209 : _GEN_177; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_242 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_210 : _GEN_178; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_243 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_211 : _GEN_179; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_244 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_212 : _GEN_180; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_245 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_213 : _GEN_181; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_246 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_214 : _GEN_182; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_247 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_215 : _GEN_183; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_248 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_216 : _GEN_184; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_249 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_217 : _GEN_185; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_250 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_218 : _GEN_186; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_251 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_219 : _GEN_187; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_252 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_220 : _GEN_188; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_253 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_221 : _GEN_189; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_254 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_222 : _GEN_190; // @[RegFile.scala 25:50]
  wire [63:0] _GEN_255 = io_wen_vec_1 & |io_rd_addr_vec_1 ? _GEN_223 : _GEN_191; // @[RegFile.scala 25:50]
  wire [63:0] _regs_dtsaddr = {{32'd0}, difftestSval}; // @[RegFile.scala 41:21 RegFile.scala 41:21]
  wire [63:0] _GEN_288 = io_rs_addr_vec_0 == difftestSaddr ? {{32'd0}, difftestSval} : _GEN_31; // @[RegFile.scala 43:46 RegFile.scala 44:29 RegFile.scala 22:23]
  wire [63:0] _GEN_289 = io_rs_addr_vec_1 == difftestSaddr ? {{32'd0}, difftestSval} : _GEN_63; // @[RegFile.scala 43:46 RegFile.scala 44:29 RegFile.scala 22:23]
  wire [63:0] _GEN_290 = io_rs_addr_vec_2 == difftestSaddr ? {{32'd0}, difftestSval} : _GEN_95; // @[RegFile.scala 43:46 RegFile.scala 44:29 RegFile.scala 22:23]
  wire [63:0] _GEN_291 = io_rs_addr_vec_3 == difftestSaddr ? {{32'd0}, difftestSval} : _GEN_127; // @[RegFile.scala 43:46 RegFile.scala 44:29 RegFile.scala 22:23]
  wire [63:0] _WIRE_0 = regs_0; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_1 = regs_1; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_2 = regs_2; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_3 = regs_3; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_4 = regs_4; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_5 = regs_5; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_6 = regs_6; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_7 = regs_7; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_8 = regs_8; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_9 = regs_9; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_10 = regs_10; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_11 = regs_11; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_12 = regs_12; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_13 = regs_13; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_14 = regs_14; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_15 = regs_15; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_16 = regs_16; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_17 = regs_17; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_18 = regs_18; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_19 = regs_19; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_20 = regs_20; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_21 = regs_21; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_22 = regs_22; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_23 = regs_23; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_24 = regs_24; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_25 = regs_25; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_26 = regs_26; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_27 = regs_27; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_28 = regs_28; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_29 = regs_29; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_30 = regs_30; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  wire [63:0] _WIRE_31 = regs_31; // @[RegFile.scala 31:34 RegFile.scala 31:34]
  assign io_rs_data_vec_0 = difftestSync ? _GEN_288 : _GEN_31; // @[RegFile.scala 40:19 RegFile.scala 22:23]
  assign io_rs_data_vec_1 = difftestSync ? _GEN_289 : _GEN_63; // @[RegFile.scala 40:19 RegFile.scala 22:23]
  assign io_rs_data_vec_2 = difftestSync ? _GEN_290 : _GEN_95; // @[RegFile.scala 40:19 RegFile.scala 22:23]
  assign io_rs_data_vec_3 = difftestSync ? _GEN_291 : _GEN_127; // @[RegFile.scala 40:19 RegFile.scala 22:23]
  assign _WIRE_0_0 = _GEN_0;
  assign _WIRE_0_1 = _WIRE_1;
  assign _WIRE_0_2 = _WIRE_2;
  assign _WIRE_0_3 = _WIRE_3;
  assign _WIRE_0_4 = _WIRE_4;
  assign _WIRE_0_5 = _WIRE_5;
  assign _WIRE_0_6 = _WIRE_6;
  assign _WIRE_0_7 = _WIRE_7;
  assign _WIRE_0_8 = _WIRE_8;
  assign _WIRE_0_9 = _WIRE_9;
  assign _WIRE_0_10 = _WIRE_10;
  assign _WIRE_0_11 = _WIRE_11;
  assign _WIRE_0_12 = _WIRE_12;
  assign _WIRE_0_13 = _WIRE_13;
  assign _WIRE_0_14 = _WIRE_14;
  assign _WIRE_0_15 = _WIRE_15;
  assign _WIRE_0_16 = _WIRE_16;
  assign _WIRE_0_17 = _WIRE_17;
  assign _WIRE_0_18 = _WIRE_18;
  assign _WIRE_0_19 = _WIRE_19;
  assign _WIRE_0_20 = _WIRE_20;
  assign _WIRE_0_21 = _WIRE_21;
  assign _WIRE_0_22 = _WIRE_22;
  assign _WIRE_0_23 = _WIRE_23;
  assign _WIRE_0_24 = _WIRE_24;
  assign _WIRE_0_25 = _WIRE_25;
  assign _WIRE_0_26 = _WIRE_26;
  assign _WIRE_0_27 = _WIRE_27;
  assign _WIRE_0_28 = _WIRE_28;
  assign _WIRE_0_29 = _WIRE_29;
  assign _WIRE_0_30 = _WIRE_30;
  assign _WIRE_0_31 = _WIRE_31;
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 20:21]
      regs_0 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h0 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_0 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_0 <= _GEN_224;
      end
    end else begin
      regs_0 <= _GEN_224;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_1 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_1 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_1 <= _GEN_225;
      end
    end else begin
      regs_1 <= _GEN_225;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_2 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h2 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_2 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_2 <= _GEN_226;
      end
    end else begin
      regs_2 <= _GEN_226;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_3 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h3 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_3 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_3 <= _GEN_227;
      end
    end else begin
      regs_3 <= _GEN_227;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_4 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h4 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_4 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_4 <= _GEN_228;
      end
    end else begin
      regs_4 <= _GEN_228;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_5 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h5 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_5 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_5 <= _GEN_229;
      end
    end else begin
      regs_5 <= _GEN_229;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_6 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h6 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_6 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_6 <= _GEN_230;
      end
    end else begin
      regs_6 <= _GEN_230;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_7 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h7 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_7 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_7 <= _GEN_231;
      end
    end else begin
      regs_7 <= _GEN_231;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_8 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h8 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_8 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_8 <= _GEN_232;
      end
    end else begin
      regs_8 <= _GEN_232;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_9 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h9 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_9 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_9 <= _GEN_233;
      end
    end else begin
      regs_9 <= _GEN_233;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_10 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'ha == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_10 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_10 <= _GEN_234;
      end
    end else begin
      regs_10 <= _GEN_234;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_11 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'hb == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_11 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_11 <= _GEN_235;
      end
    end else begin
      regs_11 <= _GEN_235;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_12 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'hc == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_12 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_12 <= _GEN_236;
      end
    end else begin
      regs_12 <= _GEN_236;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_13 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'hd == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_13 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_13 <= _GEN_237;
      end
    end else begin
      regs_13 <= _GEN_237;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_14 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'he == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_14 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_14 <= _GEN_238;
      end
    end else begin
      regs_14 <= _GEN_238;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_15 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'hf == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_15 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_15 <= _GEN_239;
      end
    end else begin
      regs_15 <= _GEN_239;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_16 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h10 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_16 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_16 <= _GEN_240;
      end
    end else begin
      regs_16 <= _GEN_240;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_17 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h11 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_17 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_17 <= _GEN_241;
      end
    end else begin
      regs_17 <= _GEN_241;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_18 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h12 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_18 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_18 <= _GEN_242;
      end
    end else begin
      regs_18 <= _GEN_242;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_19 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h13 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_19 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_19 <= _GEN_243;
      end
    end else begin
      regs_19 <= _GEN_243;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_20 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h14 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_20 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_20 <= _GEN_244;
      end
    end else begin
      regs_20 <= _GEN_244;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_21 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h15 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_21 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_21 <= _GEN_245;
      end
    end else begin
      regs_21 <= _GEN_245;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_22 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h16 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_22 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_22 <= _GEN_246;
      end
    end else begin
      regs_22 <= _GEN_246;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_23 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h17 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_23 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_23 <= _GEN_247;
      end
    end else begin
      regs_23 <= _GEN_247;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_24 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h18 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_24 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_24 <= _GEN_248;
      end
    end else begin
      regs_24 <= _GEN_248;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_25 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h19 == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_25 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_25 <= _GEN_249;
      end
    end else begin
      regs_25 <= _GEN_249;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_26 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1a == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_26 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_26 <= _GEN_250;
      end
    end else begin
      regs_26 <= _GEN_250;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_27 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1b == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_27 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_27 <= _GEN_251;
      end
    end else begin
      regs_27 <= _GEN_251;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_28 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1c == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_28 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_28 <= _GEN_252;
      end
    end else begin
      regs_28 <= _GEN_252;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_29 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1d == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_29 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_29 <= _GEN_253;
      end
    end else begin
      regs_29 <= _GEN_253;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_30 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1e == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_30 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_30 <= _GEN_254;
      end
    end else begin
      regs_30 <= _GEN_254;
    end
    if (reset) begin // @[RegFile.scala 20:21]
      regs_31 <= 64'h0; // @[RegFile.scala 20:21]
    end else if (difftestSync) begin // @[RegFile.scala 40:19]
      if (5'h1f == difftestSaddr) begin // @[RegFile.scala 41:21]
        regs_31 <= _regs_dtsaddr; // @[RegFile.scala 41:21]
      end else begin
        regs_31 <= _GEN_255;
      end
    end else begin
      regs_31 <= _GEN_255;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [63:0] io_common_io_in,
  input         io_common_io_wen,
  input  [11:0] io_common_io_num,
  output [63:0] io_common_io_out,
  input         io_event_io_exception_vec_2,
  input         io_event_io_exception_vec_3,
  input         io_event_io_exception_vec_4,
  input         io_event_io_exception_vec_6,
  input         io_event_io_deal_with_int,
  input         io_event_io_is_mret,
  input         io_event_io_is_sret,
  input         io_event_io_is_ecall,
  input  [63:0] io_event_io_bad_address,
  input  [63:0] io_event_io_epc,
  output        io_event_io_call_for_int,
  output        io_event_io_except_kill,
  output [63:0] io_event_io_redirect_pc,
  output [63:0] csrs_0_mstatus,
  output [63:0] csrs_0_sstatus,
  output [63:0] csrs_0_mepc,
  output [63:0] csrs_0_sepc,
  output [63:0] csrs_0_mtval,
  output [63:0] csrs_0_stval,
  output [63:0] csrs_0_mtvec,
  output [63:0] csrs_0_stvec,
  output [63:0] csrs_0_mcause,
  output [63:0] csrs_0_scause,
  output [63:0] csrs_0_satp,
  output [63:0] csrs_0_mip,
  output [63:0] csrs_0_mie,
  output [63:0] csrs_0_mscratch,
  output [63:0] csrs_0_sscratch,
  output [63:0] csrs_0_mideleg,
  output [63:0] csrs_0_medeleg,
  output [1:0]  current_mode_0,
  output        REG_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] current_mode; // @[CSR.scala 96:29]
  wire  true_deal_with_int = io_event_io_deal_with_int & io_event_io_call_for_int; // @[CSR.scala 97:54]
  reg [63:0] mstatus; // @[CSR.scala 113:27]
  reg [63:0] medeleg; // @[CSR.scala 114:23]
  reg [63:0] mideleg; // @[CSR.scala 115:23]
  reg [63:0] mie; // @[CSR.scala 116:27]
  reg [63:0] mtvec; // @[CSR.scala 117:23]
  reg [63:0] mcounteren; // @[CSR.scala 118:27]
  reg [63:0] mscratch; // @[CSR.scala 120:21]
  reg [63:0] mepc; // @[CSR.scala 121:21]
  reg [63:0] mcause; // @[CSR.scala 122:25]
  reg [63:0] mtval; // @[CSR.scala 123:21]
  reg [63:0] mipReg; // @[CSR.scala 125:24]
  reg [63:0] mip; // @[CSR.scala 129:24]
  reg [63:0] mcycle; // @[CSR.scala 132:30]
  reg [63:0] mcountinhibit; // @[CSR.scala 133:30]
  reg [63:0] stvec; // @[CSR.scala 140:27]
  reg [63:0] scounteren; // @[CSR.scala 141:27]
  reg [63:0] sscratch; // @[CSR.scala 143:25]
  reg [63:0] sepc; // @[CSR.scala 144:25]
  reg [63:0] scause; // @[CSR.scala 145:25]
  reg [63:0] stval; // @[CSR.scala 146:25]
  reg [63:0] satp; // @[CSR.scala 149:21]
  wire [63:0] _T_35 = 64'h222 & mideleg; // @[CSR.scala 201:50]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[CSR.scala 221:20]
  wire  _wen_T_3 = io_common_io_in[63:60] == 4'h0 | io_common_io_in[63:60] == 4'h8; // @[CSRSpec.scala 333:18]
  wire  wen = io_common_io_wen & (io_common_io_num != 12'h180 | _wen_T_3); // @[CSR.scala 228:32]
  wire [63:0] _rdata_T_2 = satp; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_3 = sscratch; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_4 = medeleg; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_5 = stvec; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_6 = sepc; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_7 = mcause; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_10 = mie & _T_35; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_11 = mipReg & _T_35; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_12 = mstatus & 64'h80000003000de122; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_13 = mtvec; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_14 = mie; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_15 = stval; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_17 = mstatus; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_20 = mideleg; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_22 = mscratch; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_25 = mepc; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_26 = mtval; // @[CSRRegMap.scala 39:84]
  wire [63:0] _rdata_T_28 = scause; // @[CSRRegMap.scala 39:84]
  wire  _rdata_T_29 = 12'hc00 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_30 = 12'hf12 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_31 = 12'h180 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_32 = 12'h140 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_33 = 12'h302 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_34 = 12'h105 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_35 = 12'h141 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_36 = 12'h342 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_37 = 12'h306 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_38 = 12'hf11 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_39 = 12'h104 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_40 = 12'h144 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_41 = 12'h100 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_42 = 12'h305 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_43 = 12'h304 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_44 = 12'h143 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_45 = 12'h301 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_46 = 12'h300 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_47 = 12'hb00 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_48 = 12'h344 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_49 = 12'h303 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_50 = 12'hf13 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_51 = 12'h340 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_52 = 12'h320 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_53 = 12'hf14 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_54 = 12'h341 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_55 = 12'h343 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_56 = 12'h106 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire  _rdata_T_57 = 12'h142 == io_common_io_num; // @[LookupTree.scala 8:34]
  wire [63:0] _rdata_T_58 = _rdata_T_29 ? mcycle : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_60 = _rdata_T_31 ? satp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_61 = _rdata_T_32 ? sscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_62 = _rdata_T_33 ? medeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_63 = _rdata_T_34 ? stvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_64 = _rdata_T_35 ? sepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_65 = _rdata_T_36 ? mcause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_66 = _rdata_T_37 ? mcounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_68 = _rdata_T_39 ? _rdata_T_10 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_69 = _rdata_T_40 ? _rdata_T_11 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_70 = _rdata_T_41 ? _rdata_T_12 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_71 = _rdata_T_42 ? mtvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_72 = _rdata_T_43 ? mie : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_73 = _rdata_T_44 ? stval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_74 = _rdata_T_45 ? 64'h800000000014112d : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_75 = _rdata_T_46 ? mstatus : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_76 = _rdata_T_47 ? mcycle : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_77 = _rdata_T_48 ? mipReg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_78 = _rdata_T_49 ? mideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_80 = _rdata_T_51 ? mscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_81 = _rdata_T_52 ? mcountinhibit : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_83 = _rdata_T_54 ? mepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_84 = _rdata_T_55 ? mtval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_85 = _rdata_T_56 ? scounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_86 = _rdata_T_57 ? scause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_88 = _rdata_T_58 | _rdata_T_60; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_89 = _rdata_T_88 | _rdata_T_61; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_90 = _rdata_T_89 | _rdata_T_62; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_91 = _rdata_T_90 | _rdata_T_63; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_92 = _rdata_T_91 | _rdata_T_64; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_93 = _rdata_T_92 | _rdata_T_65; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_94 = _rdata_T_93 | _rdata_T_66; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_96 = _rdata_T_94 | _rdata_T_68; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_97 = _rdata_T_96 | _rdata_T_69; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_98 = _rdata_T_97 | _rdata_T_70; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_99 = _rdata_T_98 | _rdata_T_71; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_100 = _rdata_T_99 | _rdata_T_72; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_101 = _rdata_T_100 | _rdata_T_73; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_102 = _rdata_T_101 | _rdata_T_74; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_103 = _rdata_T_102 | _rdata_T_75; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_104 = _rdata_T_103 | _rdata_T_76; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_105 = _rdata_T_104 | _rdata_T_77; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_106 = _rdata_T_105 | _rdata_T_78; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_108 = _rdata_T_106 | _rdata_T_80; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_109 = _rdata_T_108 | _rdata_T_81; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_111 = _rdata_T_109 | _rdata_T_83; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_112 = _rdata_T_111 | _rdata_T_84; // @[Mux.scala 27:72]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_85; // @[Mux.scala 27:72]
  wire [63:0] rdata = _rdata_T_113 | _rdata_T_86; // @[Mux.scala 27:72]
  wire [63:0] _medeleg_T = io_common_io_in & 64'hbbff; // @[CSRRegMap.scala 8:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'h4400; // @[CSRRegMap.scala 8:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[CSRRegMap.scala 8:26]
  wire [63:0] _GEN_4 = wen & io_common_io_num == 12'h141 ? io_common_io_in : sepc; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 144:25]
  wire [63:0] _GEN_5 = wen & io_common_io_num == 12'h342 ? io_common_io_in : mcause; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 122:25]
  wire [63:0] _mie_T_1 = io_common_io_in & _T_35; // @[CSRRegMap.scala 8:14]
  wire [63:0] _mie_T_2 = ~_T_35; // @[CSRRegMap.scala 8:40]
  wire [63:0] _mie_T_3 = mie & _mie_T_2; // @[CSRRegMap.scala 8:37]
  wire [63:0] _mie_T_4 = _mie_T_1 | _mie_T_3; // @[CSRRegMap.scala 8:26]
  wire [63:0] _mipReg_T_3 = mipReg & _mie_T_2; // @[CSRRegMap.scala 8:37]
  wire [63:0] _mipReg_T_4 = _mie_T_1 | _mipReg_T_3; // @[CSRRegMap.scala 8:26]
  wire [63:0] _mstatus_T_1 = io_common_io_in & 64'hc6122; // @[CSRRegMap.scala 8:14]
  wire [63:0] _mstatus_T_3 = mstatus & 64'h39edd; // @[CSRRegMap.scala 8:37]
  wire [63:0] _mstatus_T_4 = _mstatus_T_1 | _mstatus_T_3; // @[CSRRegMap.scala 8:26]
  wire [1:0] mstatus_mstatus_old_FS = _mstatus_T_4[14:13]; // @[CSRSpec.scala 206:48]
  wire  mstatus_mstatus_new_hi = mstatus_mstatus_old_FS == 2'h3; // @[CSRSpec.scala 207:42]
  wire [62:0] mstatus_mstatus_new_lo = _mstatus_T_4[62:0]; // @[CSRSpec.scala 207:62]
  wire [63:0] mstatus_mstatus_new = {mstatus_mstatus_new_hi,mstatus_mstatus_new_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_9 = wen & io_common_io_num == 12'h100 ? mstatus_mstatus_new : mstatus; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 113:27]
  wire [63:0] _GEN_12 = wen & io_common_io_num == 12'h143 ? io_common_io_in : stval; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 146:25]
  wire [1:0] mstatus_mstatus_old_1_FS = io_common_io_in[14:13]; // @[CSRSpec.scala 206:48]
  wire  mstatus_mstatus_new_hi_1 = mstatus_mstatus_old_1_FS == 2'h3; // @[CSRSpec.scala 207:42]
  wire [62:0] mstatus_mstatus_new_lo_1 = io_common_io_in[62:0]; // @[CSRSpec.scala 207:62]
  wire [63:0] mstatus_mstatus_new_1 = {mstatus_mstatus_new_hi_1,mstatus_mstatus_new_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_13 = wen & io_common_io_num == 12'h300 ? mstatus_mstatus_new_1 : _GEN_9; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11]
  wire [63:0] _mipReg_T_5 = io_common_io_in & 64'h77f; // @[CSRRegMap.scala 8:14]
  wire [63:0] _mipReg_T_7 = mipReg & 64'h80; // @[CSRRegMap.scala 8:37]
  wire [63:0] _mipReg_T_8 = _mipReg_T_5 | _mipReg_T_7; // @[CSRRegMap.scala 8:26]
  wire [63:0] _mideleg_T = io_common_io_in & 64'h222; // @[CSRRegMap.scala 8:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'h1dd; // @[CSRRegMap.scala 8:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[CSRRegMap.scala 8:26]
  wire [63:0] _GEN_18 = wen & io_common_io_num == 12'h341 ? io_common_io_in : mepc; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 121:21]
  wire [63:0] _GEN_19 = wen & io_common_io_num == 12'h343 ? io_common_io_in : mtval; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 123:21]
  wire [63:0] _GEN_21 = wen & io_common_io_num == 12'h142 ? io_common_io_in : scause; // @[CSRRegMap.scala 41:71 CSRRegMap.scala 42:11 CSR.scala 145:25]
  reg [11:0] int_cause; // @[CSR.scala 303:27]
  wire [11:0] _mip_old_MEIP_T = {{11'd0}, int_cause[11]}; // @[CSR.scala 310:50]
  wire  mip_old_MEIP = true_deal_with_int & _mip_old_MEIP_T[0]; // @[CSR.scala 310:38]
  wire [11:0] _mip_old_SEIP_T = {{9'd0}, int_cause[11:9]}; // @[CSR.scala 311:50]
  wire  mip_old_SEIP = true_deal_with_int & _mip_old_SEIP_T[0]; // @[CSR.scala 311:38]
  wire [11:0] _mip_old_MTIP_T = {{7'd0}, int_cause[11:7]}; // @[CSR.scala 313:50]
  wire  mip_old_MTIP = true_deal_with_int & _mip_old_MTIP_T[0]; // @[CSR.scala 313:38]
  wire [11:0] _mip_old_STIP_T = {{5'd0}, int_cause[11:5]}; // @[CSR.scala 314:50]
  wire  mip_old_STIP = true_deal_with_int & _mip_old_STIP_T[0]; // @[CSR.scala 314:38]
  wire [11:0] _mip_old_MSIP_T = {{3'd0}, int_cause[11:3]}; // @[CSR.scala 312:50]
  wire  mip_old_MSIP = true_deal_with_int & _mip_old_MSIP_T[0]; // @[CSR.scala 312:38]
  wire [5:0] mip_new_lo = {mip_old_STIP,1'h0,mip_old_MSIP,3'h0}; // @[CSR.scala 335:28]
  wire [63:0] _mip_new_T = {52'h0,mip_old_MEIP,1'h0,mip_old_SEIP,1'h0,mip_old_MTIP,1'h0,mip_new_lo}; // @[CSR.scala 335:28]
  wire [63:0] interrupt_deleg = mideleg & mip; // @[CSR.scala 317:33]
  wire  mip_mask_11 = ~interrupt_deleg[9]; // @[CSR.scala 328:22]
  wire  mip_mask_9 = ~mip_mask_11; // @[CSR.scala 330:22]
  wire  mip_mask_7 = ~interrupt_deleg[5]; // @[CSR.scala 328:22]
  wire  mip_mask_5 = ~mip_mask_7; // @[CSR.scala 330:22]
  wire  mip_mask_3 = ~interrupt_deleg[1]; // @[CSR.scala 328:22]
  wire  mip_mask_1 = ~mip_mask_3; // @[CSR.scala 330:22]
  wire [5:0] mip_new_lo_1 = {mip_mask_5,1'h0,mip_mask_3,1'h0,mip_mask_1,1'h0}; // @[CSR.scala 335:48]
  wire [11:0] _mip_new_T_1 = {mip_mask_11,1'h0,mip_mask_9,1'h0,mip_mask_7,1'h0,mip_new_lo_1}; // @[CSR.scala 335:48]
  wire [63:0] _GEN_54 = {{52'd0}, _mip_new_T_1}; // @[CSR.scala 335:31]
  wire [63:0] _mip_new_T_2 = _mip_new_T & _GEN_54; // @[CSR.scala 335:31]
  wire [63:0] mip_new = _mip_new_T_2 & mie; // @[CSR.scala 335:51]
  wire [63:0] mipOut = mip_new | mip; // @[CSR.scala 336:21]
  wire [63:0] _io_common_io_out_T = mipOut & 64'h222; // @[CSR.scala 235:41]
  wire [63:0] _io_common_io_out_T_2 = _rdata_T_48 ? mipOut : rdata; // @[Mux.scala 80:57]
  wire [63:0] _io_common_io_out_T_4 = _rdata_T_40 ? _io_common_io_out_T : _io_common_io_out_T_2; // @[Mux.scala 80:57]
  wire  old_mstatus_UIE = mstatus[0]; // @[CSR.scala 245:51]
  wire  old_mstatus_SIE = mstatus[1]; // @[CSR.scala 245:51]
  wire  old_mstatus_WPRI2 = mstatus[2]; // @[CSR.scala 245:51]
  wire  old_mstatus_MIE = mstatus[3]; // @[CSR.scala 245:51]
  wire  old_mstatus_UPIE = mstatus[4]; // @[CSR.scala 245:51]
  wire  old_mstatus_SPIE = mstatus[5]; // @[CSR.scala 245:51]
  wire  old_mstatus_WPRI6 = mstatus[6]; // @[CSR.scala 245:51]
  wire  old_mstatus_MPIE = mstatus[7]; // @[CSR.scala 245:51]
  wire  old_mstatus_SPP = mstatus[8]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_WPRI9 = mstatus[10:9]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_MPP = mstatus[12:11]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_FS = mstatus[14:13]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_XS = mstatus[16:15]; // @[CSR.scala 245:51]
  wire  old_mstatus_MPRV = mstatus[17]; // @[CSR.scala 245:51]
  wire  old_mstatus_SUM = mstatus[18]; // @[CSR.scala 245:51]
  wire  old_mstatus_MXR = mstatus[19]; // @[CSR.scala 245:51]
  wire  old_mstatus_TVM = mstatus[20]; // @[CSR.scala 245:51]
  wire  old_mstatus_TW = mstatus[21]; // @[CSR.scala 245:51]
  wire  old_mstatus_TSR = mstatus[22]; // @[CSR.scala 245:51]
  wire [8:0] old_mstatus_WPRI23 = mstatus[31:23]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_UXL = mstatus[33:32]; // @[CSR.scala 245:51]
  wire [1:0] old_mstatus_SXL = mstatus[35:34]; // @[CSR.scala 245:51]
  wire [26:0] old_mstatus_WPRI36 = mstatus[62:36]; // @[CSR.scala 245:51]
  wire  old_mstatus_SD = mstatus[63]; // @[CSR.scala 245:51]
  wire [5:0] mstatus_lo_lo_1 = {old_mstatus_SPIE,old_mstatus_UPIE,old_mstatus_MPIE,old_mstatus_WPRI2,old_mstatus_SIE,
    old_mstatus_UIE}; // @[CSR.scala 251:34]
  wire [14:0] mstatus_lo_1 = {old_mstatus_FS,2'h0,old_mstatus_WPRI9,old_mstatus_SPP,1'h1,old_mstatus_WPRI6,
    mstatus_lo_lo_1}; // @[CSR.scala 251:34]
  wire [6:0] mstatus_hi_lo_1 = {old_mstatus_TW,old_mstatus_TVM,old_mstatus_MXR,old_mstatus_SUM,old_mstatus_MPRV,
    old_mstatus_XS}; // @[CSR.scala 251:34]
  wire [63:0] _mstatus_T_9 = {old_mstatus_SD,old_mstatus_WPRI36,old_mstatus_SXL,old_mstatus_UXL,old_mstatus_WPRI23,
    old_mstatus_TSR,mstatus_hi_lo_1,mstatus_lo_1}; // @[CSR.scala 251:34]
  wire [63:0] _GEN_24 = io_event_io_is_mret ? mepc : 64'h0; // @[CSR.scala 244:29 CSR.scala 252:16]
  wire [1:0] _current_mode_T = {1'h0,old_mstatus_SPP}; // @[Cat.scala 30:58]
  wire [5:0] mstatus_lo_lo_2 = {1'h1,old_mstatus_UPIE,old_mstatus_MIE,old_mstatus_WPRI2,old_mstatus_SPIE,old_mstatus_UIE
    }; // @[CSR.scala 263:36]
  wire [14:0] mstatus_lo_2 = {old_mstatus_FS,old_mstatus_MPP,old_mstatus_WPRI9,1'h0,old_mstatus_MPIE,old_mstatus_WPRI6,
    mstatus_lo_lo_2}; // @[CSR.scala 263:36]
  wire [63:0] _mstatus_T_10 = {old_mstatus_SD,old_mstatus_WPRI36,old_mstatus_SXL,old_mstatus_UXL,old_mstatus_WPRI23,
    old_mstatus_TSR,mstatus_hi_lo_1,mstatus_lo_2}; // @[CSR.scala 263:36]
  wire [63:0] ret_target = io_event_io_is_sret ? sepc : _GEN_24; // @[CSR.scala 256:31 CSR.scala 264:18]
  wire  _illegal_csr_num_illegalAddr_T_1 = _rdata_T_29 ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_3 = _rdata_T_30 ? 1'h0 : _illegal_csr_num_illegalAddr_T_1; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_5 = _rdata_T_31 ? 1'h0 : _illegal_csr_num_illegalAddr_T_3; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_7 = _rdata_T_32 ? 1'h0 : _illegal_csr_num_illegalAddr_T_5; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_9 = _rdata_T_33 ? 1'h0 : _illegal_csr_num_illegalAddr_T_7; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_11 = _rdata_T_34 ? 1'h0 : _illegal_csr_num_illegalAddr_T_9; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_13 = _rdata_T_35 ? 1'h0 : _illegal_csr_num_illegalAddr_T_11; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_15 = _rdata_T_36 ? 1'h0 : _illegal_csr_num_illegalAddr_T_13; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_17 = _rdata_T_37 ? 1'h0 : _illegal_csr_num_illegalAddr_T_15; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_19 = _rdata_T_38 ? 1'h0 : _illegal_csr_num_illegalAddr_T_17; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_21 = _rdata_T_39 ? 1'h0 : _illegal_csr_num_illegalAddr_T_19; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_23 = _rdata_T_40 ? 1'h0 : _illegal_csr_num_illegalAddr_T_21; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_25 = _rdata_T_41 ? 1'h0 : _illegal_csr_num_illegalAddr_T_23; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_27 = _rdata_T_42 ? 1'h0 : _illegal_csr_num_illegalAddr_T_25; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_29 = _rdata_T_43 ? 1'h0 : _illegal_csr_num_illegalAddr_T_27; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_31 = _rdata_T_44 ? 1'h0 : _illegal_csr_num_illegalAddr_T_29; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_33 = _rdata_T_45 ? 1'h0 : _illegal_csr_num_illegalAddr_T_31; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_35 = _rdata_T_46 ? 1'h0 : _illegal_csr_num_illegalAddr_T_33; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_37 = _rdata_T_47 ? 1'h0 : _illegal_csr_num_illegalAddr_T_35; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_39 = _rdata_T_48 ? 1'h0 : _illegal_csr_num_illegalAddr_T_37; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_41 = _rdata_T_49 ? 1'h0 : _illegal_csr_num_illegalAddr_T_39; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_43 = _rdata_T_50 ? 1'h0 : _illegal_csr_num_illegalAddr_T_41; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_45 = _rdata_T_51 ? 1'h0 : _illegal_csr_num_illegalAddr_T_43; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_47 = _rdata_T_52 ? 1'h0 : _illegal_csr_num_illegalAddr_T_45; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_49 = _rdata_T_53 ? 1'h0 : _illegal_csr_num_illegalAddr_T_47; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_51 = _rdata_T_54 ? 1'h0 : _illegal_csr_num_illegalAddr_T_49; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_53 = _rdata_T_55 ? 1'h0 : _illegal_csr_num_illegalAddr_T_51; // @[Mux.scala 80:57]
  wire  _illegal_csr_num_illegalAddr_T_55 = _rdata_T_56 ? 1'h0 : _illegal_csr_num_illegalAddr_T_53; // @[Mux.scala 80:57]
  wire  illegal_csr_num_illegalAddr = _rdata_T_57 ? 1'h0 : _illegal_csr_num_illegalAddr_T_55; // @[Mux.scala 80:57]
  wire  illegal_csr_num = illegal_csr_num_illegalAddr & io_common_io_wen; // @[CSR.scala 283:76]
  wire  _csrExcpVec_11_T = current_mode == 2'h3; // @[CSR.scala 291:53]
  wire  csrExcpVec_11 = current_mode == 2'h3 & io_event_io_is_ecall; // @[CSR.scala 291:69]
  wire  _csrExcpVec_9_T = current_mode == 2'h1; // @[CSR.scala 292:53]
  wire  csrExcpVec_9 = current_mode == 2'h1 & io_event_io_is_ecall; // @[CSR.scala 292:69]
  wire  csrExcpVec_8 = current_mode == 2'h0 & io_event_io_is_ecall; // @[CSR.scala 293:69]
  wire [15:0] _allExcpVec_T = {4'h0,csrExcpVec_11,1'h0,csrExcpVec_9,csrExcpVec_8,4'h0,1'h0,illegal_csr_num,2'h0}; // @[CSR.scala 297:42]
  wire [15:0] _allExcpVec_T_1 = {8'h0,1'h0,io_event_io_exception_vec_6,1'h0,io_event_io_exception_vec_4,
    io_event_io_exception_vec_3,io_event_io_exception_vec_2,2'h0}; // @[CSR.scala 297:69]
  wire [15:0] allExcpVec = _allExcpVec_T | _allExcpVec_T_1; // @[CSR.scala 297:45]
  wire  has_excp = |allExcpVec; // @[CSR.scala 298:39]
  wire [2:0] _excp_no_T_1 = allExcpVec[5] ? 3'h5 : 3'h0; // @[CSR.scala 299:93]
  wire [2:0] _excp_no_T_3 = allExcpVec[7] ? 3'h7 : _excp_no_T_1; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_5 = allExcpVec[13] ? 4'hd : {{1'd0}, _excp_no_T_3}; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_7 = allExcpVec[15] ? 4'hf : _excp_no_T_5; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_9 = allExcpVec[4] ? 4'h4 : _excp_no_T_7; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_11 = allExcpVec[6] ? 4'h6 : _excp_no_T_9; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_13 = allExcpVec[11] ? 4'hb : _excp_no_T_11; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_15 = allExcpVec[9] ? 4'h9 : _excp_no_T_13; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_17 = allExcpVec[8] ? 4'h8 : _excp_no_T_15; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_19 = allExcpVec[0] ? 4'h0 : _excp_no_T_17; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_21 = allExcpVec[2] ? 4'h2 : _excp_no_T_19; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_23 = allExcpVec[1] ? 4'h1 : _excp_no_T_21; // @[CSR.scala 299:93]
  wire [3:0] _excp_no_T_25 = allExcpVec[12] ? 4'hc : _excp_no_T_23; // @[CSR.scala 299:93]
  wire [3:0] excp_no = allExcpVec[3] ? 4'h3 : _excp_no_T_25; // @[CSR.scala 299:93]
  wire  detect_int_5 = mip[5]; // @[CSR.scala 306:51]
  wire [5:0] int_cause_lo = {detect_int_5,1'h0,1'h0,3'h0}; // @[CSR.scala 303:39]
  wire [11:0] _int_cause_T = {6'h0,detect_int_5,1'h0,1'h0,3'h0}; // @[CSR.scala 303:39]
  wire [63:0] mipWire = mip_new & 64'hfffffffffffffdff; // @[CSR.scala 337:22]
  wire [63:0] _mip_T = mipWire | mipReg; // @[CSR.scala 338:19]
  wire [5:0] mip_lo = {_mip_T[5],_mip_T[4],_mip_T[3],_mip_T[2],_mip_T[1],_mip_T[0]}; // @[CSR.scala 338:59]
  wire [63:0] _mip_T_14 = {_mip_T[63:12],_mip_T[11],_mip_T[10],_mip_T[9],_mip_T[8],_mip_T[7],_mip_T[6],mip_lo}; // @[CSR.scala 338:59]
  wire  _intrVecEnable_0_T_56 = current_mode < 2'h3; // @[CSR.scala 341:107]
  wire  _intrVecEnable_0_T_57 = _csrExcpVec_11_T & old_mstatus_MIE | current_mode < 2'h3; // @[CSR.scala 341:90]
  wire  intrVecEnable_0 = interrupt_deleg[0] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_1 = interrupt_deleg[1] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_2 = interrupt_deleg[2] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_3 = interrupt_deleg[3] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_4 = interrupt_deleg[4] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_5 = interrupt_deleg[5] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_6 = interrupt_deleg[6] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_7 = interrupt_deleg[7] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_8 = interrupt_deleg[8] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_9 = interrupt_deleg[9] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_10 = interrupt_deleg[10] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire  intrVecEnable_11 = interrupt_deleg[11] ? _csrExcpVec_9_T & old_mstatus_SIE | current_mode < 2'h1 :
    _intrVecEnable_0_T_57; // @[CSR.scala 340:40]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _int_cause_T; // @[CSR.scala 345:28]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[CSR.scala 345:70]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[CSR.scala 345:70]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[CSR.scala 345:48]
  wire  has_intr = |intrVec; // @[CSR.scala 347:38]
  wire [11:0] _intr_no_T = {{5'd0}, intrVec[11:5]}; // @[CSR.scala 348:100]
  wire [3:0] _intr_no_T_2 = _intr_no_T[0] ? 4'h5 : 4'h0; // @[CSR.scala 348:92]
  wire [11:0] _intr_no_T_3 = {{1'd0}, intrVec[11:1]}; // @[CSR.scala 348:100]
  wire [3:0] _intr_no_T_5 = _intr_no_T_3[0] ? 4'h1 : _intr_no_T_2; // @[CSR.scala 348:92]
  wire [11:0] _intr_no_T_6 = {{9'd0}, intrVec[11:9]}; // @[CSR.scala 348:100]
  wire [3:0] _intr_no_T_8 = _intr_no_T_6[0] ? 4'h9 : _intr_no_T_5; // @[CSR.scala 348:92]
  wire [11:0] _intr_no_T_9 = {{7'd0}, intrVec[11:7]}; // @[CSR.scala 348:100]
  wire [3:0] _intr_no_T_11 = _intr_no_T_9[0] ? 4'h7 : _intr_no_T_8; // @[CSR.scala 348:92]
  wire [11:0] _intr_no_T_12 = {{3'd0}, intrVec[11:3]}; // @[CSR.scala 348:100]
  wire [3:0] _intr_no_T_14 = _intr_no_T_12[0] ? 4'h3 : _intr_no_T_11; // @[CSR.scala 348:92]
  wire [11:0] _intr_no_T_15 = {{11'd0}, intrVec[11]}; // @[CSR.scala 348:100]
  wire [3:0] intr_no = _intr_no_T_15[0] ? 4'hb : _intr_no_T_14; // @[CSR.scala 348:92]
  wire  has_excp_intr = has_excp | has_intr; // @[CSR.scala 352:32]
  wire [3:0] _cause_no_T = has_intr ? intr_no : excp_no; // @[CSR.scala 354:18]
  wire [63:0] _deleg_to_s_T = has_intr ? mideleg : medeleg; // @[CSR.scala 355:23]
  wire [63:0] cause_no = {{60'd0}, _cause_no_T}; // @[CSR.scala 353:27 CSR.scala 354:12]
  wire [63:0] _deleg_to_s_T_2 = _deleg_to_s_T >> cause_no[3:0]; // @[CSR.scala 355:51]
  wire  deleg_to_s = _deleg_to_s_T_2[0] & _intrVecEnable_0_T_56; // @[CSR.scala 355:68]
  wire  _T_106 = true_deal_with_int | has_excp; // @[CSR.scala 357:27]
  wire [63:0] _tval_T_1 = 64'hc == cause_no ? io_event_io_bad_address : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_3 = 64'hd == cause_no ? io_event_io_bad_address : _tval_T_1; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_5 = 64'hf == cause_no ? io_event_io_bad_address : _tval_T_3; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_7 = 64'h0 == cause_no ? io_event_io_bad_address : _tval_T_5; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_9 = 64'h4 == cause_no ? io_event_io_bad_address : _tval_T_7; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_11 = 64'h6 == cause_no ? io_event_io_bad_address : _tval_T_9; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_13 = 64'h1 == cause_no ? io_event_io_bad_address : _tval_T_11; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_15 = 64'h5 == cause_no ? io_event_io_bad_address : _tval_T_13; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_17 = 64'h7 == cause_no ? io_event_io_bad_address : _tval_T_15; // @[Mux.scala 80:57]
  wire [63:0] _tval_T_19 = 64'h3 == cause_no ? io_event_io_bad_address : _tval_T_17; // @[Mux.scala 80:57]
  wire [63:0] tval = 64'h2 == cause_no ? 64'h0 : _tval_T_19; // @[Mux.scala 80:57]
  wire [62:0] scause_lo = cause_no[62:0]; // @[CSR.scala 384:39]
  wire [63:0] _scause_T_5 = {has_intr,scause_lo}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_29 = deleg_to_s ? current_mode : {{1'd0}, old_mstatus_SPP}; // @[CSR.scala 383:22 CSR.scala 385:23]
  wire  new_mstatus_2_SPIE = deleg_to_s ? old_mstatus_SIE : old_mstatus_SPIE; // @[CSR.scala 383:22 CSR.scala 386:24]
  wire  new_mstatus_2_SIE = deleg_to_s ? 1'h0 : old_mstatus_SIE; // @[CSR.scala 383:22 CSR.scala 387:23]
  wire [1:0] new_mstatus_2_MPP = deleg_to_s ? old_mstatus_MPP : current_mode; // @[CSR.scala 383:22 CSR.scala 393:23]
  wire  new_mstatus_2_MPIE = deleg_to_s ? old_mstatus_MPIE : old_mstatus_MIE; // @[CSR.scala 383:22 CSR.scala 394:24]
  wire  new_mstatus_2_MIE = deleg_to_s & old_mstatus_MIE; // @[CSR.scala 383:22 CSR.scala 395:23]
  wire [5:0] mstatus_lo_lo_3 = {new_mstatus_2_SPIE,old_mstatus_UPIE,new_mstatus_2_MIE,old_mstatus_WPRI2,
    new_mstatus_2_SIE,old_mstatus_UIE}; // @[CSR.scala 400:34]
  wire  new_mstatus_2_SPP = _GEN_29[0];
  wire [14:0] mstatus_lo_3 = {old_mstatus_FS,new_mstatus_2_MPP,old_mstatus_WPRI9,new_mstatus_2_SPP,new_mstatus_2_MPIE,
    old_mstatus_WPRI6,mstatus_lo_lo_3}; // @[CSR.scala 400:34]
  wire [63:0] _mstatus_T_11 = {old_mstatus_SD,old_mstatus_WPRI36,old_mstatus_SXL,old_mstatus_UXL,old_mstatus_WPRI23,
    old_mstatus_TSR,mstatus_hi_lo_1,mstatus_lo_3}; // @[CSR.scala 400:34]
  wire [63:0] tvec = deleg_to_s ? stvec : mtvec; // @[CSR.scala 404:24]
  wire [2:0] _trap_target_T_2 = {tvec[0], 2'h0}; // @[CSR.scala 405:63]
  wire [66:0] _trap_target_T_3 = _trap_target_T_2 * cause_no; // @[CSR.scala 405:69]
  wire [66:0] _trap_target_T_5 = 67'hfffffffffffffffc + _trap_target_T_3; // @[CSR.scala 405:43]
  wire [66:0] _GEN_61 = {{3'd0}, tvec}; // @[CSR.scala 405:26]
  wire [66:0] trap_target = _GEN_61 & _trap_target_T_5; // @[CSR.scala 405:26]
  wire [66:0] _io_event_io_redirect_pc_T = has_excp_intr ? trap_target : {{3'd0}, ret_target}; // @[CSR.scala 406:33]
  reg  REG; // @[CSR.scala 413:34]
  wire [63:0] _csrs_sstatus_T_70 = _rdata_T_12; // @[CSRRegMap.scala 53:75]
  wire [63:0] csrs_mstatus = mstatus; // @[CSR.scala 417:20 CSR.scala 418:19]
  wire [63:0] csrs_sstatus = _rdata_T_12; // @[CSRRegMap.scala 53:75]
  wire [63:0] csrs_mepc = mepc; // @[CSR.scala 417:20 CSR.scala 420:19]
  wire [63:0] csrs_sepc = sepc; // @[CSR.scala 417:20 CSR.scala 421:19]
  wire [63:0] csrs_mtval = mtval; // @[CSR.scala 417:20 CSR.scala 422:19]
  wire [63:0] csrs_stval = stval; // @[CSR.scala 417:20 CSR.scala 423:19]
  wire [63:0] csrs_mtvec = mtvec; // @[CSR.scala 417:20 CSR.scala 424:19]
  wire [63:0] csrs_stvec = stvec; // @[CSR.scala 417:20 CSR.scala 425:19]
  wire [63:0] csrs_mcause = mcause; // @[CSR.scala 417:20 CSR.scala 426:19]
  wire [63:0] csrs_scause = scause; // @[CSR.scala 417:20 CSR.scala 427:19]
  wire [63:0] csrs_satp = satp; // @[CSR.scala 417:20 CSR.scala 428:19]
  wire [63:0] csrs_mip = mip; // @[CSR.scala 417:20 CSR.scala 429:19]
  wire [63:0] csrs_mie = mie; // @[CSR.scala 417:20 CSR.scala 430:19]
  wire [63:0] csrs_mscratch = mscratch; // @[CSR.scala 417:20 CSR.scala 431:19]
  wire [63:0] csrs_sscratch = sscratch; // @[CSR.scala 417:20 CSR.scala 432:19]
  wire [63:0] csrs_mideleg = mideleg; // @[CSR.scala 417:20 CSR.scala 433:19]
  wire [63:0] csrs_medeleg = medeleg; // @[CSR.scala 417:20 CSR.scala 434:19]
  assign io_common_io_out = _rdata_T_47 ? 64'h1 : _io_common_io_out_T_4; // @[Mux.scala 80:57]
  assign io_event_io_call_for_int = |intrVec; // @[CSR.scala 347:38]
  assign io_event_io_except_kill = _T_106 | io_event_io_is_mret | io_event_io_is_sret; // @[CSR.scala 407:84]
  assign io_event_io_redirect_pc = _io_event_io_redirect_pc_T[63:0]; // @[CSR.scala 406:27]
  assign csrs_0_mstatus = _rdata_T_17;
  assign csrs_0_sstatus = _csrs_sstatus_T_70;
  assign csrs_0_mepc = _rdata_T_25;
  assign csrs_0_sepc = _rdata_T_6;
  assign csrs_0_mtval = _rdata_T_26;
  assign csrs_0_stval = _rdata_T_15;
  assign csrs_0_mtvec = _rdata_T_13;
  assign csrs_0_stvec = _rdata_T_5;
  assign csrs_0_mcause = _rdata_T_7;
  assign csrs_0_scause = _rdata_T_28;
  assign csrs_0_satp = _rdata_T_2;
  assign csrs_0_mip = mip;
  assign csrs_0_mie = _rdata_T_14;
  assign csrs_0_mscratch = _rdata_T_22;
  assign csrs_0_sscratch = _rdata_T_3;
  assign csrs_0_mideleg = _rdata_T_20;
  assign csrs_0_medeleg = _rdata_T_4;
  assign current_mode_0 = current_mode;
  assign REG_0 = REG;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 96:29]
      current_mode <= 2'h3; // @[CSR.scala 96:29]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        current_mode <= 2'h1; // @[CSR.scala 389:20]
      end else begin
        current_mode <= 2'h3; // @[CSR.scala 397:20]
      end
    end else if (io_event_io_is_sret) begin // @[CSR.scala 256:31]
      current_mode <= _current_mode_T; // @[CSR.scala 262:20]
    end else if (io_event_io_is_mret) begin // @[CSR.scala 244:29]
      current_mode <= old_mstatus_MPP; // @[CSR.scala 250:18]
    end
    if (reset) begin // @[CSR.scala 113:27]
      mstatus <= 64'h0; // @[CSR.scala 113:27]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      mstatus <= _mstatus_T_11; // @[CSR.scala 400:13]
    end else if (io_event_io_is_sret) begin // @[CSR.scala 256:31]
      mstatus <= _mstatus_T_10; // @[CSR.scala 263:15]
    end else if (io_event_io_is_mret) begin // @[CSR.scala 244:29]
      mstatus <= _mstatus_T_9; // @[CSR.scala 251:13]
    end else begin
      mstatus <= _GEN_13;
    end
    if (wen & io_common_io_num == 12'h302) begin // @[CSRRegMap.scala 41:71]
      medeleg <= _medeleg_T_3; // @[CSRRegMap.scala 42:11]
    end
    if (wen & io_common_io_num == 12'h303) begin // @[CSRRegMap.scala 41:71]
      mideleg <= _mideleg_T_3; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 116:27]
      mie <= 64'h0; // @[CSR.scala 116:27]
    end else if (wen & io_common_io_num == 12'h304) begin // @[CSRRegMap.scala 41:71]
      mie <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end else if (wen & io_common_io_num == 12'h104) begin // @[CSRRegMap.scala 41:71]
      mie <= _mie_T_4; // @[CSRRegMap.scala 42:11]
    end
    if (wen & io_common_io_num == 12'h305) begin // @[CSRRegMap.scala 41:71]
      mtvec <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 118:27]
      mcounteren <= 64'h0; // @[CSR.scala 118:27]
    end else if (wen & io_common_io_num == 12'h306) begin // @[CSRRegMap.scala 41:71]
      mcounteren <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (wen & io_common_io_num == 12'h340) begin // @[CSRRegMap.scala 41:71]
      mscratch <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        mepc <= _GEN_18;
      end else begin
        mepc <= io_event_io_epc; // @[CSR.scala 396:12]
      end
    end else begin
      mepc <= _GEN_18;
    end
    if (reset) begin // @[CSR.scala 122:25]
      mcause <= 64'h0; // @[CSR.scala 122:25]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        mcause <= _GEN_5;
      end else begin
        mcause <= _scause_T_5; // @[CSR.scala 392:14]
      end
    end else begin
      mcause <= _GEN_5;
    end
    if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        mtval <= _GEN_19;
      end else if (true_deal_with_int) begin // @[CSR.scala 390:19]
        mtval <= 64'h0;
      end else if (64'h2 == cause_no) begin // @[Mux.scala 80:57]
        mtval <= 64'h0;
      end else begin
        mtval <= _tval_T_19;
      end
    end else begin
      mtval <= _GEN_19;
    end
    if (reset) begin // @[CSR.scala 125:24]
      mipReg <= 64'h0; // @[CSR.scala 125:24]
    end else if (wen & io_common_io_num == 12'h344) begin // @[CSRRegMap.scala 41:71]
      mipReg <= _mipReg_T_8; // @[CSRRegMap.scala 42:11]
    end else if (wen & io_common_io_num == 12'h144) begin // @[CSRRegMap.scala 41:71]
      mipReg <= _mipReg_T_4; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 129:24]
      mip <= 64'h0; // @[CSR.scala 129:24]
    end else begin
      mip <= _mip_T_14; // @[CSR.scala 338:7]
    end
    if (reset) begin // @[CSR.scala 132:30]
      mcycle <= 64'h0; // @[CSR.scala 132:30]
    end else begin
      mcycle <= _mcycle_T_1; // @[CSR.scala 221:10]
    end
    if (reset) begin // @[CSR.scala 133:30]
      mcountinhibit <= 64'h0; // @[CSR.scala 133:30]
    end else if (wen & io_common_io_num == 12'h320) begin // @[CSRRegMap.scala 41:71]
      mcountinhibit <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 140:27]
      stvec <= 64'h0; // @[CSR.scala 140:27]
    end else if (wen & io_common_io_num == 12'h105) begin // @[CSRRegMap.scala 41:71]
      stvec <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 141:27]
      scounteren <= 64'h0; // @[CSR.scala 141:27]
    end else if (wen & io_common_io_num == 12'h106) begin // @[CSRRegMap.scala 41:71]
      scounteren <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 143:25]
      sscratch <= 64'h0; // @[CSR.scala 143:25]
    end else if (wen & io_common_io_num == 12'h140) begin // @[CSRRegMap.scala 41:71]
      sscratch <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    if (reset) begin // @[CSR.scala 144:25]
      sepc <= 64'h0; // @[CSR.scala 144:25]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        sepc <= io_event_io_epc; // @[CSR.scala 388:12]
      end else begin
        sepc <= _GEN_4;
      end
    end else begin
      sepc <= _GEN_4;
    end
    if (reset) begin // @[CSR.scala 145:25]
      scause <= 64'h0; // @[CSR.scala 145:25]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        scause <= _scause_T_5; // @[CSR.scala 384:14]
      end else begin
        scause <= _GEN_21;
      end
    end else begin
      scause <= _GEN_21;
    end
    if (reset) begin // @[CSR.scala 146:25]
      stval <= 64'h0; // @[CSR.scala 146:25]
    end else if (true_deal_with_int | has_excp) begin // @[CSR.scala 357:40]
      if (deleg_to_s) begin // @[CSR.scala 383:22]
        if (true_deal_with_int) begin // @[CSR.scala 390:19]
          stval <= 64'h0;
        end else begin
          stval <= tval;
        end
      end else begin
        stval <= _GEN_12;
      end
    end else begin
      stval <= _GEN_12;
    end
    if (reset) begin // @[CSR.scala 149:21]
      satp <= 64'h0; // @[CSR.scala 149:21]
    end else if (wen & io_common_io_num == 12'h180) begin // @[CSRRegMap.scala 41:71]
      satp <= io_common_io_in; // @[CSRRegMap.scala 42:11]
    end
    int_cause <= {6'h0,int_cause_lo}; // @[CSR.scala 303:39]
    REG <= io_event_io_deal_with_int & io_event_io_call_for_int; // @[CSR.scala 97:54]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  current_mode = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mstatus = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  medeleg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mideleg = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mie = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mtvec = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcounteren = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mscratch = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mepc = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mcause = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mtval = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mipReg = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  mip = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mcycle = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  mcountinhibit = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  stvec = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  scounteren = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  sscratch = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  sepc = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  scause = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stval = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  int_cause = _RAND_22[11:0];
  _RAND_23 = {1{`RANDOM}};
  REG = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Backend(
  input          clock,
  input          reset,
  output         io_fb_bmfs_redirect_kill,
  output [31:0]  io_fb_bmfs_redirect_pc,
  output         io_fb_bmfs_bpu_v,
  output         io_fb_bmfs_bpu_errpr,
  output [63:0]  io_fb_bmfs_bpu_pc_br,
  output [63:0]  io_fb_bmfs_bpu_target,
  output         io_fb_bmfs_bpu_taken,
  input  [1:0]   io_fb_fmbs_instn,
  input  [160:0] io_fb_fmbs_inst_ops_0,
  input  [160:0] io_fb_fmbs_inst_ops_1,
  output         io_fb_fmbs_please_wait,
  output         io_dcache_req_valid,
  output [31:0]  io_dcache_req_bits_addr,
  output [63:0]  io_dcache_req_bits_wdata,
  output         io_dcache_req_bits_wen,
  output [2:0]   io_dcache_req_bits_mtype,
  input          io_dcache_resp_valid,
  input  [31:0]  io_dcache_resp_bits_rdata_0,
  input  [31:0]  io_dcache_resp_bits_rdata_1,
  output [63:0]  csrs_mstatus,
  output [63:0]  csrs_sstatus,
  output [63:0]  csrs_mepc,
  output [63:0]  csrs_sepc,
  output [63:0]  csrs_mtval,
  output [63:0]  csrs_stval,
  output [63:0]  csrs_mtvec,
  output [63:0]  csrs_stvec,
  output [63:0]  csrs_mcause,
  output [63:0]  csrs_scause,
  output [63:0]  csrs_satp,
  output [63:0]  csrs_mip,
  output [63:0]  csrs_mie,
  output [63:0]  csrs_mscratch,
  output [63:0]  csrs_sscratch,
  output [63:0]  csrs_mideleg,
  output [63:0]  csrs_medeleg,
  output [63:0]  istall_0,
  output         _WIRE_4_0_0,
  output         _WIRE_4_0_1,
  output         _WIRE_4_0_2,
  output [31:0]  _WIRE_1_0_0,
  output [31:0]  _WIRE_1_0_1,
  output [31:0]  _WIRE_1_0_2,
  input  [4:0]   difftest_saddr,
  output [1:0]   current_mode,
  output [63:0]  _WIRE_0_0,
  output [63:0]  _WIRE_0_1,
  output [63:0]  _WIRE_0_2,
  output [63:0]  _WIRE_0_3,
  output [63:0]  _WIRE_0_4,
  output [63:0]  _WIRE_0_5,
  output [63:0]  _WIRE_0_6,
  output [63:0]  _WIRE_0_7,
  output [63:0]  _WIRE_0_8,
  output [63:0]  _WIRE_0_9,
  output [63:0]  _WIRE_0_10,
  output [63:0]  _WIRE_0_11,
  output [63:0]  _WIRE_0_12,
  output [63:0]  _WIRE_0_13,
  output [63:0]  _WIRE_0_14,
  output [63:0]  _WIRE_0_15,
  output [63:0]  _WIRE_0_16,
  output [63:0]  _WIRE_0_17,
  output [63:0]  _WIRE_0_18,
  output [63:0]  _WIRE_0_19,
  output [63:0]  _WIRE_0_20,
  output [63:0]  _WIRE_0_21,
  output [63:0]  _WIRE_0_22,
  output [63:0]  _WIRE_0_23,
  output [63:0]  _WIRE_0_24,
  output [63:0]  _WIRE_0_25,
  output [63:0]  _WIRE_0_26,
  output [63:0]  _WIRE_0_27,
  output [63:0]  _WIRE_0_28,
  output [63:0]  _WIRE_0_29,
  output [63:0]  _WIRE_0_30,
  output [63:0]  _WIRE_0_31,
  output [63:0]  dstall_0,
  output         _WIRE_6_0,
  output         _WIRE_6_1,
  output         _WIRE_6_2,
  output [63:0]  counter_0,
  input          icache_stall,
  input  [31:0]  difftest_sval,
  output [63:0]  mduStall_0,
  output [31:0]  _WIRE_3_0_0,
  output [31:0]  _WIRE_3_0_1,
  output [31:0]  _WIRE_3_0_2,
  output [63:0]  common_0,
  output         _WIRE_5_0_0,
  output         _WIRE_5_0_1,
  output         _WIRE_5_0_2,
  output [63:0]  instret_0,
  output [1:0]   _WIRE_2_0_0,
  output [1:0]   _WIRE_2_0_1,
  output [1:0]   _WIRE_2_0_2,
  output         REG_0,
  input          difftest_sync,
  output         wbInsts_0_ysyx_debug
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] alu_io_a; // @[Backend.scala 59:28]
  wire [63:0] alu_io_b; // @[Backend.scala 59:28]
  wire [4:0] alu_io_aluOp; // @[Backend.scala 59:28]
  wire  alu_io_aluExpand; // @[Backend.scala 59:28]
  wire  alu_io_aluCsr; // @[Backend.scala 59:28]
  wire [63:0] alu_io_csr; // @[Backend.scala 59:28]
  wire [63:0] alu_io_r; // @[Backend.scala 59:28]
  wire  alu_io_zero; // @[Backend.scala 59:28]
  wire  mdu_clock; // @[Backend.scala 60:28]
  wire  mdu_reset; // @[Backend.scala 60:28]
  wire  mdu_io_kill; // @[Backend.scala 60:28]
  wire  mdu_io_req_valid; // @[Backend.scala 60:28]
  wire [4:0] mdu_io_req_op; // @[Backend.scala 60:28]
  wire  mdu_io_req_expand; // @[Backend.scala 60:28]
  wire [63:0] mdu_io_req_in1; // @[Backend.scala 60:28]
  wire [63:0] mdu_io_req_in2; // @[Backend.scala 60:28]
  wire [63:0] mdu_io_resp_r; // @[Backend.scala 60:28]
  wire  mdu_io_resp_valid; // @[Backend.scala 60:28]
  wire  issueQueue_clock; // @[Backend.scala 68:28]
  wire  issueQueue_reset; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_illegal; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_dout_0_next_pc; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_0_alu_mdu_lsu; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_dout_0_branch_type; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_0_src_a; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_0_src_b; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_write_dest; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_0_alu_op; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_alu_expand; // @[Backend.scala 68:28]
  wire [2:0] issueQueue_io_dout_0_mem_width; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_0_write_src; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_0_rs1; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_0_rs2; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_0_rd; // @[Backend.scala 68:28]
  wire [19:0] issueQueue_io_dout_0_imm; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_0_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_predict_taken; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_0_target_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_ysyx_debug; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_0_ysyx_print; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_0_inst; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_illegal; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_dout_1_next_pc; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_1_alu_mdu_lsu; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_dout_1_branch_type; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_1_src_a; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_1_src_b; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_write_dest; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_1_alu_op; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_alu_expand; // @[Backend.scala 68:28]
  wire [2:0] issueQueue_io_dout_1_mem_width; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_dout_1_write_src; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_1_rs1; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_1_rs2; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_dout_1_rd; // @[Backend.scala 68:28]
  wire [19:0] issueQueue_io_dout_1_imm; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_1_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_predict_taken; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_1_target_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_ysyx_debug; // @[Backend.scala 68:28]
  wire  issueQueue_io_dout_1_ysyx_print; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_dout_1_inst; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_enqStep; // @[Backend.scala 68:28]
  wire  issueQueue_io_enqReq; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_deqStep; // @[Backend.scala 68:28]
  wire  issueQueue_io_deqReq; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_illegal; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_din_0_next_pc; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_0_alu_mdu_lsu; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_din_0_branch_type; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_0_src_a; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_0_src_b; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_write_dest; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_0_alu_op; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_alu_expand; // @[Backend.scala 68:28]
  wire [2:0] issueQueue_io_din_0_mem_width; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_0_write_src; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_0_rs1; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_0_rs2; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_0_rd; // @[Backend.scala 68:28]
  wire [19:0] issueQueue_io_din_0_imm; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_0_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_predict_taken; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_0_target_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_ysyx_debug; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_0_ysyx_print; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_0_inst; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_illegal; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_din_1_next_pc; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_1_alu_mdu_lsu; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_din_1_branch_type; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_1_src_a; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_1_src_b; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_write_dest; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_1_alu_op; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_alu_expand; // @[Backend.scala 68:28]
  wire [2:0] issueQueue_io_din_1_mem_width; // @[Backend.scala 68:28]
  wire [1:0] issueQueue_io_din_1_write_src; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_1_rs1; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_1_rs2; // @[Backend.scala 68:28]
  wire [4:0] issueQueue_io_din_1_rd; // @[Backend.scala 68:28]
  wire [19:0] issueQueue_io_din_1_imm; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_1_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_predict_taken; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_1_target_pc; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_ysyx_debug; // @[Backend.scala 68:28]
  wire  issueQueue_io_din_1_ysyx_print; // @[Backend.scala 68:28]
  wire [31:0] issueQueue_io_din_1_inst; // @[Backend.scala 68:28]
  wire  issueQueue_io_flush; // @[Backend.scala 68:28]
  wire  issueQueue_io_sufficient; // @[Backend.scala 68:28]
  wire [3:0] issueQueue_io_items; // @[Backend.scala 68:28]
  wire  issueArbiter_io_insts_in_0_illegal; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_in_0_next_pc; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_0_alu_mdu_lsu; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_in_0_branch_type; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_0_src_a; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_0_src_b; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_0_write_dest; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_0_alu_op; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_0_alu_expand; // @[Backend.scala 69:28]
  wire [2:0] issueArbiter_io_insts_in_0_mem_width; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_0_write_src; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_0_rs1; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_0_rs2; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_0_rd; // @[Backend.scala 69:28]
  wire [19:0] issueArbiter_io_insts_in_0_imm; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_0_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_0_predict_taken; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_0_target_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_0_ysyx_debug; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_0_ysyx_print; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_0_inst; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_illegal; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_in_1_next_pc; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_1_alu_mdu_lsu; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_in_1_branch_type; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_1_src_a; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_1_src_b; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_write_dest; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_1_alu_op; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_alu_expand; // @[Backend.scala 69:28]
  wire [2:0] issueArbiter_io_insts_in_1_mem_width; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_in_1_write_src; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_1_rs1; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_1_rs2; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_in_1_rd; // @[Backend.scala 69:28]
  wire [19:0] issueArbiter_io_insts_in_1_imm; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_1_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_predict_taken; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_1_target_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_ysyx_debug; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_in_1_ysyx_print; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_in_1_inst; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_queue_items; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_ld_dest_ex; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rss_in_0; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rss_in_1; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rts_in_0; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rts_in_1; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rss_out_0; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rss_out_1; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rss_out_2; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rts_out_0; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rts_out_1; // @[Backend.scala 69:28]
  wire [63:0] issueArbiter_io_rts_out_2; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_illegal; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_out_0_next_pc; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_0_alu_mdu_lsu; // @[Backend.scala 69:28]
  wire [3:0] issueArbiter_io_insts_out_0_branch_type; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_0_src_a; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_0_src_b; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_write_dest; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_0_alu_op; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_alu_expand; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_0_write_src; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_0_rs1; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_0_rd; // @[Backend.scala 69:28]
  wire [19:0] issueArbiter_io_insts_out_0_imm; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_0_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_predict_taken; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_0_target_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_ysyx_debug; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_0_ysyx_print; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_0_inst; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_1_src_a; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_1_src_b; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_1_write_dest; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_1_alu_op; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_1_alu_expand; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_1_rd; // @[Backend.scala 69:28]
  wire [19:0] issueArbiter_io_insts_out_1_imm; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_1_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_1_ysyx_print; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_1_inst; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_out_2_src_a; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_2_write_dest; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_2_alu_op; // @[Backend.scala 69:28]
  wire [2:0] issueArbiter_io_insts_out_2_mem_width; // @[Backend.scala 69:28]
  wire [4:0] issueArbiter_io_insts_out_2_rd; // @[Backend.scala 69:28]
  wire [19:0] issueArbiter_io_insts_out_2_imm; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_2_pc; // @[Backend.scala 69:28]
  wire  issueArbiter_io_insts_out_2_ysyx_print; // @[Backend.scala 69:28]
  wire [31:0] issueArbiter_io_insts_out_2_inst; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_issue_num; // @[Backend.scala 69:28]
  wire  issueArbiter_io_issue_fu_valid_0; // @[Backend.scala 69:28]
  wire  issueArbiter_io_issue_fu_valid_1; // @[Backend.scala 69:28]
  wire  issueArbiter_io_issue_fu_valid_2; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_order_0; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_order_1; // @[Backend.scala 69:28]
  wire [1:0] issueArbiter_io_insts_order_2; // @[Backend.scala 69:28]
  wire  regFile_clock; // @[Backend.scala 131:32]
  wire  regFile_reset; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rs_addr_vec_0; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rs_addr_vec_1; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rs_addr_vec_2; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rs_addr_vec_3; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rs_data_vec_0; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rs_data_vec_1; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rs_data_vec_2; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rs_data_vec_3; // @[Backend.scala 131:32]
  wire  regFile_io_wen_vec_0; // @[Backend.scala 131:32]
  wire  regFile_io_wen_vec_1; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rd_addr_vec_0; // @[Backend.scala 131:32]
  wire [4:0] regFile_io_rd_addr_vec_1; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rd_data_vec_0; // @[Backend.scala 131:32]
  wire [63:0] regFile_io_rd_data_vec_1; // @[Backend.scala 131:32]
  wire [4:0] regFile_difftestSaddr; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_0; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_1; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_2; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_3; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_4; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_5; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_6; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_7; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_8; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_9; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_10; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_11; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_12; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_13; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_14; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_15; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_16; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_17; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_18; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_19; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_20; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_21; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_22; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_23; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_24; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_25; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_26; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_27; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_28; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_29; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_30; // @[Backend.scala 131:32]
  wire [63:0] regFile__WIRE_0_31; // @[Backend.scala 131:32]
  wire [31:0] regFile_difftestSval; // @[Backend.scala 131:32]
  wire  regFile_difftestSync; // @[Backend.scala 131:32]
  wire  csr_clock; // @[Backend.scala 132:32]
  wire  csr_reset; // @[Backend.scala 132:32]
  wire [63:0] csr_io_common_io_in; // @[Backend.scala 132:32]
  wire  csr_io_common_io_wen; // @[Backend.scala 132:32]
  wire [11:0] csr_io_common_io_num; // @[Backend.scala 132:32]
  wire [63:0] csr_io_common_io_out; // @[Backend.scala 132:32]
  wire  csr_io_event_io_exception_vec_2; // @[Backend.scala 132:32]
  wire  csr_io_event_io_exception_vec_3; // @[Backend.scala 132:32]
  wire  csr_io_event_io_exception_vec_4; // @[Backend.scala 132:32]
  wire  csr_io_event_io_exception_vec_6; // @[Backend.scala 132:32]
  wire  csr_io_event_io_deal_with_int; // @[Backend.scala 132:32]
  wire  csr_io_event_io_is_mret; // @[Backend.scala 132:32]
  wire  csr_io_event_io_is_sret; // @[Backend.scala 132:32]
  wire  csr_io_event_io_is_ecall; // @[Backend.scala 132:32]
  wire [63:0] csr_io_event_io_bad_address; // @[Backend.scala 132:32]
  wire [63:0] csr_io_event_io_epc; // @[Backend.scala 132:32]
  wire  csr_io_event_io_call_for_int; // @[Backend.scala 132:32]
  wire  csr_io_event_io_except_kill; // @[Backend.scala 132:32]
  wire [63:0] csr_io_event_io_redirect_pc; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mstatus; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_sstatus; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mepc; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_sepc; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mtval; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_stval; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mtvec; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_stvec; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mcause; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_scause; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_satp; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mip; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mie; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mscratch; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_sscratch; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_mideleg; // @[Backend.scala 132:32]
  wire [63:0] csr_csrs_0_medeleg; // @[Backend.scala 132:32]
  wire [1:0] csr_current_mode_0; // @[Backend.scala 132:32]
  wire  csr_REG_0; // @[Backend.scala 132:32]
  reg  exInsts_0_illegal; // @[Backend.scala 81:29]
  reg [3:0] exInsts_0_next_pc; // @[Backend.scala 81:29]
  reg [1:0] exInsts_0_alu_mdu_lsu; // @[Backend.scala 81:29]
  reg [3:0] exInsts_0_branch_type; // @[Backend.scala 81:29]
  reg [1:0] exInsts_0_src_a; // @[Backend.scala 81:29]
  reg [1:0] exInsts_0_src_b; // @[Backend.scala 81:29]
  reg  exInsts_0_write_dest; // @[Backend.scala 81:29]
  reg [4:0] exInsts_0_alu_op; // @[Backend.scala 81:29]
  reg  exInsts_0_alu_expand; // @[Backend.scala 81:29]
  reg [1:0] exInsts_0_write_src; // @[Backend.scala 81:29]
  reg [4:0] exInsts_0_rs1; // @[Backend.scala 81:29]
  reg [4:0] exInsts_0_rd; // @[Backend.scala 81:29]
  reg [19:0] exInsts_0_imm; // @[Backend.scala 81:29]
  reg [31:0] exInsts_0_pc; // @[Backend.scala 81:29]
  reg  exInsts_0_predict_taken; // @[Backend.scala 81:29]
  reg [31:0] exInsts_0_target_pc; // @[Backend.scala 81:29]
  reg  exInsts_0_ysyx_debug; // @[Backend.scala 81:29]
  reg  exInsts_0_ysyx_print; // @[Backend.scala 81:29]
  reg [31:0] exInsts_0_inst; // @[Backend.scala 81:29]
  reg [1:0] exInsts_1_src_a; // @[Backend.scala 81:29]
  reg [1:0] exInsts_1_src_b; // @[Backend.scala 81:29]
  reg  exInsts_1_write_dest; // @[Backend.scala 81:29]
  reg [4:0] exInsts_1_alu_op; // @[Backend.scala 81:29]
  reg  exInsts_1_alu_expand; // @[Backend.scala 81:29]
  reg [4:0] exInsts_1_rd; // @[Backend.scala 81:29]
  reg [19:0] exInsts_1_imm; // @[Backend.scala 81:29]
  reg [31:0] exInsts_1_pc; // @[Backend.scala 81:29]
  reg  exInsts_1_ysyx_print; // @[Backend.scala 81:29]
  reg [31:0] exInsts_1_inst; // @[Backend.scala 81:29]
  reg [1:0] exInsts_2_src_a; // @[Backend.scala 81:29]
  reg  exInsts_2_write_dest; // @[Backend.scala 81:29]
  reg [4:0] exInsts_2_alu_op; // @[Backend.scala 81:29]
  reg [2:0] exInsts_2_mem_width; // @[Backend.scala 81:29]
  reg [4:0] exInsts_2_rd; // @[Backend.scala 81:29]
  reg [19:0] exInsts_2_imm; // @[Backend.scala 81:29]
  reg [31:0] exInsts_2_pc; // @[Backend.scala 81:29]
  reg  exInsts_2_ysyx_print; // @[Backend.scala 81:29]
  reg [31:0] exInsts_2_inst; // @[Backend.scala 81:29]
  reg [1:0] exInstsOrder_0; // @[Backend.scala 82:95]
  reg [1:0] exInstsOrder_1; // @[Backend.scala 82:95]
  reg [1:0] exInstsOrder_2; // @[Backend.scala 82:95]
  reg  exInstsValid_0; // @[Backend.scala 83:29]
  reg  exInstsValid_1; // @[Backend.scala 83:29]
  reg  exInstsValid_2; // @[Backend.scala 83:29]
  reg [63:0] exFwdRsData_0; // @[Backend.scala 84:25]
  reg [63:0] exFwdRsData_1; // @[Backend.scala 84:25]
  reg [63:0] exFwdRsData_2; // @[Backend.scala 84:25]
  reg [63:0] exFwdRtData_0; // @[Backend.scala 85:25]
  reg [63:0] exFwdRtData_1; // @[Backend.scala 85:25]
  reg [63:0] exFwdRtData_2; // @[Backend.scala 85:25]
  wire  isExPCBr = exInsts_0_next_pc == 4'h2; // @[Backend.scala 86:41]
  wire  _isExPCJump_T_1 = exInsts_0_next_pc == 4'h3; // @[Backend.scala 87:87]
  wire  isExPCJump = exInsts_0_next_pc == 4'h4 | exInsts_0_next_pc == 4'h3; // @[Backend.scala 87:65]
  wire [31:0] genImm_0_hi_hi = exInsts_0_imm[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_0_T_5 = {genImm_0_hi_hi,exInsts_0_imm,12'h0}; // @[Cat.scala 30:58]
  wire [43:0] genImm_0_hi_1 = exInsts_0_imm[19] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_0_T_8 = {genImm_0_hi_1,exInsts_0_imm}; // @[Cat.scala 30:58]
  wire [63:0] genImm_0 = exInsts_0_alu_op == 5'ha | exInsts_0_src_a == 2'h2 ? _genImm_0_T_5 : _genImm_0_T_8; // @[Backend.scala 54:8]
  wire [63:0] _GEN_410 = {{32'd0}, exInsts_0_pc}; // @[Backend.scala 91:36]
  wire [63:0] brPC = _GEN_410 + genImm_0; // @[Backend.scala 91:36]
  wire  exCsrValid = exInsts_0_src_b == 2'h2; // @[Backend.scala 92:37]
  wire  _aluValid_T = ~io_fb_bmfs_redirect_kill; // @[Backend.scala 279:36]
  wire  aluValid = exInstsValid_0 & ~io_fb_bmfs_redirect_kill; // @[Backend.scala 279:33]
  wire [31:0] genImm_2_hi_hi = exInsts_2_imm[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_2_T_5 = {genImm_2_hi_hi,exInsts_2_imm,12'h0}; // @[Cat.scala 30:58]
  wire [43:0] genImm_2_hi_1 = exInsts_2_imm[19] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_2_T_8 = {genImm_2_hi_1,exInsts_2_imm}; // @[Cat.scala 30:58]
  wire [63:0] genImm_2 = exInsts_2_alu_op == 5'ha | exInsts_2_src_a == 2'h2 ? _genImm_2_T_5 : _genImm_2_T_8; // @[Backend.scala 54:8]
  wire [63:0] ldstAddr = exFwdRsData_2 + genImm_2; // @[Backend.scala 97:37]
  wire  _memMisaligned_T_9 = |ldstAddr[2:0]; // @[Backend.scala 107:46]
  wire  _memMisaligned_T_7 = |ldstAddr[1:0]; // @[Backend.scala 106:46]
  wire  _memMisaligned_T_13 = 3'h3 == exInsts_2_mem_width ? ldstAddr[0] : 3'h2 == exInsts_2_mem_width & ldstAddr[0]; // @[Mux.scala 80:57]
  wire  _memMisaligned_T_15 = 3'h4 == exInsts_2_mem_width ? _memMisaligned_T_7 : _memMisaligned_T_13; // @[Mux.scala 80:57]
  wire  _memMisaligned_T_17 = 3'h6 == exInsts_2_mem_width ? _memMisaligned_T_7 : _memMisaligned_T_15; // @[Mux.scala 80:57]
  wire  memMisaligned = 3'h5 == exInsts_2_mem_width ? _memMisaligned_T_9 : _memMisaligned_T_17; // @[Mux.scala 80:57]
  wire  _aluExptMask_T = exInstsValid_2 & memMisaligned; // @[Backend.scala 113:42]
  wire  aluExptMask = exInstsValid_2 & memMisaligned & exInstsOrder_2 < exInstsOrder_0; // @[Backend.scala 113:59]
  wire  exInstsTrueValid_0 = aluValid & ~aluExptMask; // @[Backend.scala 414:35]
  wire  _reBranchBrTaken_T_9 = ~alu_io_r[0]; // @[Backend.scala 377:44]
  wire  _reBranchBrTaken_T_5 = $signed(alu_io_r) < 64'sh0; // @[Backend.scala 375:48]
  wire  _reBranchBrTaken_T_3 = $signed(alu_io_r) >= 64'sh0; // @[Backend.scala 374:48]
  wire  _reBranchBrTaken_T_1 = ~alu_io_zero; // @[Backend.scala 373:44]
  wire  _reBranchBrTaken_T = alu_io_zero; // @[Backend.scala 371:72]
  wire  _reBranchBrTaken_T_11 = 4'h2 == exInsts_0_branch_type ? _reBranchBrTaken_T_1 : _reBranchBrTaken_T; // @[Mux.scala 80:57]
  wire  _reBranchBrTaken_T_13 = 4'h3 == exInsts_0_branch_type ? _reBranchBrTaken_T_3 : _reBranchBrTaken_T_11; // @[Mux.scala 80:57]
  wire  _reBranchBrTaken_T_15 = 4'h6 == exInsts_0_branch_type ? _reBranchBrTaken_T_5 : _reBranchBrTaken_T_13; // @[Mux.scala 80:57]
  wire  _reBranchBrTaken_T_17 = 4'h4 == exInsts_0_branch_type ? alu_io_r[0] : _reBranchBrTaken_T_15; // @[Mux.scala 80:57]
  wire  _reBranchBrTaken_T_19 = 4'h5 == exInsts_0_branch_type ? _reBranchBrTaken_T_9 : _reBranchBrTaken_T_17; // @[Mux.scala 80:57]
  wire  _GEN_219 = isExPCBr & _reBranchBrTaken_T_19; // @[Backend.scala 370:21 Backend.scala 371:23 Backend.scala 363:19]
  wire  reBranchBrTaken = exInstsTrueValid_0 & _GEN_219; // @[Backend.scala 369:29 Backend.scala 363:19]
  wire [31:0] _exReBranchPC_T_3 = exInsts_0_pc + 32'h4; // @[Backend.scala 93:96]
  wire [63:0] _exReBranchPC_T_4 = ~reBranchBrTaken | exCsrValid ? {{32'd0}, _exReBranchPC_T_3} : brPC; // @[Backend.scala 93:49]
  wire [62:0] jumpPc_hi = genImm_0[62:0]; // @[Backend.scala 366:34]
  wire [63:0] _jumpPc_T_1 = {jumpPc_hi,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _jumpPc_T_3 = _GEN_410 + _jumpPc_T_1; // @[Backend.scala 366:19]
  wire [63:0] _jumpPc_T_5 = exFwdRsData_0 + genImm_0; // @[Backend.scala 367:25]
  wire [62:0] jumpPc_hi_1 = _jumpPc_T_5[63:1]; // @[Backend.scala 367:37]
  wire [63:0] _jumpPc_T_6 = {jumpPc_hi_1,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _jumpPc_T_7 = _isExPCJump_T_1 ? _jumpPc_T_3 : _jumpPc_T_6; // @[Backend.scala 364:16]
  wire [31:0] jumpPc = _jumpPc_T_7[31:0]; // @[Backend.scala 90:26 Backend.scala 364:10]
  wire [63:0] exReBranchPC = isExPCJump ? {{32'd0}, jumpPc} : _exReBranchPC_T_4; // @[Backend.scala 93:25]
  reg  exInterruptd; // @[Backend.scala 99:29]
  wire  mduExptMask = _aluExptMask_T & exInstsOrder_2 < exInstsOrder_1; // @[Backend.scala 114:59]
  wire  ldstValid = exInstsValid_2 & _aluValid_T; // @[Backend.scala 281:33]
  wire  exMemRealValid = ldstValid & ~memMisaligned; // @[Backend.scala 115:44]
  wire  bpuV = (isExPCBr | isExPCJump) & exInstsValid_0; // @[Backend.scala 116:44]
  wire  _bpuErrpr_T_2 = exInsts_0_target_pc[31:2] != brPC[31:2]; // @[Backend.scala 117:69]
  wire  _bpuErrpr_T_7 = exInsts_0_target_pc[31:2] != jumpPc[31:2]; // @[Backend.scala 118:71]
  wire  _bpuErrpr_T_8 = isExPCJump & exInsts_0_target_pc[31:2] != jumpPc[31:2]; // @[Backend.scala 118:30]
  reg [31:0] reBranchPC; // @[Backend.scala 124:29]
  reg [63:0] wbResult_0; // @[Backend.scala 125:29]
  reg [63:0] wbResult_1; // @[Backend.scala 125:29]
  reg  wbInstsValid_0; // @[Backend.scala 126:33]
  reg  wbInstsValid_1; // @[Backend.scala 126:33]
  reg  wbInstsValid_2; // @[Backend.scala 126:33]
  reg [1:0] wbInstsOrder_0; // @[Backend.scala 127:29]
  reg [1:0] wbInstsOrder_1; // @[Backend.scala 127:29]
  reg [1:0] wbInstsOrder_2; // @[Backend.scala 127:29]
  reg  wbInsts__0_illegal; // @[Backend.scala 128:33]
  reg [3:0] wbInsts__0_next_pc; // @[Backend.scala 128:33]
  reg [1:0] wbInsts__0_alu_mdu_lsu; // @[Backend.scala 128:33]
  reg  wbInsts__0_write_dest; // @[Backend.scala 128:33]
  reg [4:0] wbInsts__0_rd; // @[Backend.scala 128:33]
  reg [19:0] wbInsts__0_imm; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__0_pc; // @[Backend.scala 128:33]
  reg  wbInsts__0_ysyx_debug; // @[Backend.scala 128:33]
  reg  wbInsts__0_ysyx_print; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__0_inst; // @[Backend.scala 128:33]
  reg  wbInsts__1_write_dest; // @[Backend.scala 128:33]
  reg [4:0] wbInsts__1_rd; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__1_pc; // @[Backend.scala 128:33]
  reg  wbInsts__1_ysyx_print; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__1_inst; // @[Backend.scala 128:33]
  reg  wbInsts__2_write_dest; // @[Backend.scala 128:33]
  reg [2:0] wbInsts__2_mem_width; // @[Backend.scala 128:33]
  reg [4:0] wbInsts__2_rd; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__2_pc; // @[Backend.scala 128:33]
  reg  wbInsts__2_ysyx_print; // @[Backend.scala 128:33]
  reg [31:0] wbInsts__2_inst; // @[Backend.scala 128:33]
  reg  wbReBranch; // @[Backend.scala 134:33]
  reg [31:0] wbMisalignedAddr; // @[Backend.scala 137:33]
  reg  wbInterruptd; // @[Backend.scala 138:33]
  reg  wbLdMa; // @[Backend.scala 139:33]
  reg  wbStMa; // @[Backend.scala 140:33]
  reg  wbBpuV; // @[Backend.scala 141:33]
  reg  wbBpuErrpr; // @[Backend.scala 142:33]
  wire [29:0] wbBpuPCBr_hi = exInsts_0_pc[31:2]; // @[Backend.scala 144:45]
  wire [1:0] wbBpuPCBr_lo = exInsts_0_target_pc[1:0]; // @[Backend.scala 144:84]
  reg [31:0] wbBpuPCBr; // @[Backend.scala 144:33]
  reg [63:0] wbBpuTarget; // @[Backend.scala 145:33]
  reg  wbBpuTaken; // @[Backend.scala 146:33]
  reg [63:0] wbCsrData; // @[Backend.scala 148:29]
  reg  wbMemReqValid; // @[Backend.scala 306:30]
  wire  dcacheStall = wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
  wire  _stall_i_T = ~mdu_io_resp_valid; // @[Backend.scala 359:29]
  wire  bubble_w = dcacheStall | ~mdu_io_resp_valid; // @[Backend.scala 359:26]
  wire  _issueQueue_io_deqReq_T = ~bubble_w; // @[Backend.scala 156:28]
  wire [1:0] issueNum = issueArbiter_io_issue_num; // @[Backend.scala 64:26 Backend.scala 171:31]
  wire [4:0] _issueArbiter_io_ld_dest_ex_T_1 = exInstsValid_2 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] issueInsts_0_rs1 = issueQueue_io_dout_0_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  wire [63:0] rsData_0 = regFile_io_rs_data_vec_0; // @[Backend.scala 74:26 Backend.scala 227:15]
  wire [63:0] _GEN_0 = wbInsts__0_rd == issueInsts_0_rs1 ? wbResult_0 : rsData_0; // @[Backend.scala 185:51 Backend.scala 186:24 Backend.scala 178:18]
  wire [4:0] issueInsts_0_rs2 = issueQueue_io_dout_0_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  wire [63:0] rtData_0 = regFile_io_rs_data_vec_1; // @[Backend.scala 75:26 Backend.scala 228:15]
  wire [63:0] _GEN_1 = wbInsts__0_rd == issueInsts_0_rs2 ? wbResult_0 : rtData_0; // @[Backend.scala 188:51 Backend.scala 189:24 Backend.scala 179:18]
  wire [4:0] issueInsts_1_rs1 = issueQueue_io_dout_1_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  wire [63:0] rsData_1 = regFile_io_rs_data_vec_2; // @[Backend.scala 74:26 Backend.scala 227:15]
  wire [63:0] _GEN_2 = wbInsts__0_rd == issueInsts_1_rs1 ? wbResult_0 : rsData_1; // @[Backend.scala 185:51 Backend.scala 186:24 Backend.scala 178:18]
  wire [4:0] issueInsts_1_rs2 = issueQueue_io_dout_1_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  wire [63:0] rtData_1 = regFile_io_rs_data_vec_3; // @[Backend.scala 75:26 Backend.scala 228:15]
  wire [63:0] _GEN_3 = wbInsts__0_rd == issueInsts_1_rs2 ? wbResult_0 : rtData_1; // @[Backend.scala 188:51 Backend.scala 189:24 Backend.scala 179:18]
  wire [63:0] _GEN_4 = wbInstsValid_0 & wbInsts__0_write_dest & wbInsts__0_rd != 5'h0 ? _GEN_0 : rsData_0; // @[Backend.scala 183:98 Backend.scala 178:18]
  wire [63:0] _GEN_5 = wbInstsValid_0 & wbInsts__0_write_dest & wbInsts__0_rd != 5'h0 ? _GEN_1 : rtData_0; // @[Backend.scala 183:98 Backend.scala 179:18]
  wire [63:0] _GEN_6 = wbInstsValid_0 & wbInsts__0_write_dest & wbInsts__0_rd != 5'h0 ? _GEN_2 : rsData_1; // @[Backend.scala 183:98 Backend.scala 178:18]
  wire [63:0] _GEN_7 = wbInstsValid_0 & wbInsts__0_write_dest & wbInsts__0_rd != 5'h0 ? _GEN_3 : rtData_1; // @[Backend.scala 183:98 Backend.scala 179:18]
  wire  _T_9 = wbInstsValid_1 & wbInsts__1_write_dest; // @[Backend.scala 183:26]
  wire [63:0] _GEN_8 = wbInsts__1_rd == issueInsts_0_rs1 ? wbResult_1 : _GEN_4; // @[Backend.scala 185:51 Backend.scala 186:24]
  wire [63:0] _GEN_9 = wbInsts__1_rd == issueInsts_0_rs2 ? wbResult_1 : _GEN_5; // @[Backend.scala 188:51 Backend.scala 189:24]
  wire [63:0] _GEN_10 = wbInsts__1_rd == issueInsts_1_rs1 ? wbResult_1 : _GEN_6; // @[Backend.scala 185:51 Backend.scala 186:24]
  wire [63:0] _GEN_11 = wbInsts__1_rd == issueInsts_1_rs2 ? wbResult_1 : _GEN_7; // @[Backend.scala 188:51 Backend.scala 189:24]
  wire [63:0] _GEN_12 = wbInstsValid_1 & wbInsts__1_write_dest & wbInsts__1_rd != 5'h0 ? _GEN_8 : _GEN_4; // @[Backend.scala 183:98]
  wire [63:0] _GEN_13 = wbInstsValid_1 & wbInsts__1_write_dest & wbInsts__1_rd != 5'h0 ? _GEN_9 : _GEN_5; // @[Backend.scala 183:98]
  wire [63:0] _GEN_14 = wbInstsValid_1 & wbInsts__1_write_dest & wbInsts__1_rd != 5'h0 ? _GEN_10 : _GEN_6; // @[Backend.scala 183:98]
  wire [63:0] _GEN_15 = wbInstsValid_1 & wbInsts__1_write_dest & wbInsts__1_rd != 5'h0 ? _GEN_11 : _GEN_7; // @[Backend.scala 183:98]
  wire  _T_43 = 3'h0 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [63:0] _dataFromDcache_T = {io_dcache_resp_bits_rdata_1,io_dcache_resp_bits_rdata_0}; // @[Backend.scala 439:56]
  reg [31:0] wbMemReq_addr; // @[Backend.scala 315:25]
  wire [5:0] delayed_req_bits = {wbMemReq_addr[2:0], 3'h0}; // @[Backend.scala 438:61]
  wire [63:0] dataFromDcache = _dataFromDcache_T >> delayed_req_bits; // @[Backend.scala 439:59]
  wire [55:0] wbLdData_hi = dataFromDcache[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] wbLdData_lo = dataFromDcache[7:0]; // @[Backend.scala 444:99]
  wire [63:0] _wbLdData_T_2 = {wbLdData_hi,wbLdData_lo}; // @[Cat.scala 30:58]
  wire  _T_44 = 3'h1 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [63:0] _wbLdData_T_3 = {56'h0,wbLdData_lo}; // @[Cat.scala 30:58]
  wire  _T_45 = 3'h2 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [47:0] wbLdData_hi_2 = dataFromDcache[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] wbLdData_lo_2 = dataFromDcache[15:0]; // @[Backend.scala 446:101]
  wire [63:0] _wbLdData_T_6 = {wbLdData_hi_2,wbLdData_lo_2}; // @[Cat.scala 30:58]
  wire  _T_46 = 3'h3 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [63:0] _wbLdData_T_7 = {48'h0,wbLdData_lo_2}; // @[Cat.scala 30:58]
  wire  _T_47 = 3'h4 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [31:0] wbLdData_hi_4 = dataFromDcache[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] wbLdData_lo_4 = dataFromDcache[31:0]; // @[Backend.scala 448:101]
  wire [63:0] _wbLdData_T_10 = {wbLdData_hi_4,wbLdData_lo_4}; // @[Cat.scala 30:58]
  wire  _T_48 = 3'h6 == wbInsts__2_mem_width; // @[Conditional.scala 37:30]
  wire [63:0] _wbLdData_T_11 = {32'h0,wbLdData_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_223 = _T_48 ? _wbLdData_T_11 : dataFromDcache; // @[Conditional.scala 39:67 Backend.scala 449:41 Backend.scala 442:12]
  wire [63:0] _GEN_224 = _T_47 ? _wbLdData_T_10 : _GEN_223; // @[Conditional.scala 39:67 Backend.scala 448:41]
  wire [63:0] _GEN_225 = _T_46 ? _wbLdData_T_7 : _GEN_224; // @[Conditional.scala 39:67 Backend.scala 447:41]
  wire [63:0] _GEN_226 = _T_45 ? _wbLdData_T_6 : _GEN_225; // @[Conditional.scala 39:67 Backend.scala 446:41]
  wire [63:0] _GEN_227 = _T_44 ? _wbLdData_T_3 : _GEN_226; // @[Conditional.scala 39:67 Backend.scala 445:41]
  wire [63:0] wbLdData = _T_43 ? _wbLdData_T_2 : _GEN_227; // @[Conditional.scala 40:58 Backend.scala 444:41]
  wire [63:0] _GEN_16 = wbInsts__2_rd == issueInsts_0_rs1 ? wbLdData : _GEN_12; // @[Backend.scala 185:51 Backend.scala 186:24]
  wire [63:0] _GEN_17 = wbInsts__2_rd == issueInsts_0_rs2 ? wbLdData : _GEN_13; // @[Backend.scala 188:51 Backend.scala 189:24]
  wire [63:0] _GEN_18 = wbInsts__2_rd == issueInsts_1_rs1 ? wbLdData : _GEN_14; // @[Backend.scala 185:51 Backend.scala 186:24]
  wire [63:0] _GEN_19 = wbInsts__2_rd == issueInsts_1_rs2 ? wbLdData : _GEN_15; // @[Backend.scala 188:51 Backend.scala 189:24]
  wire [63:0] _GEN_20 = wbInstsValid_2 & wbInsts__2_write_dest & wbInsts__2_rd != 5'h0 ? _GEN_16 : _GEN_12; // @[Backend.scala 183:98]
  wire [63:0] _GEN_21 = wbInstsValid_2 & wbInsts__2_write_dest & wbInsts__2_rd != 5'h0 ? _GEN_17 : _GEN_13; // @[Backend.scala 183:98]
  wire [63:0] _GEN_22 = wbInstsValid_2 & wbInsts__2_write_dest & wbInsts__2_rd != 5'h0 ? _GEN_18 : _GEN_14; // @[Backend.scala 183:98]
  wire [63:0] _GEN_23 = wbInstsValid_2 & wbInsts__2_write_dest & wbInsts__2_rd != 5'h0 ? _GEN_19 : _GEN_15; // @[Backend.scala 183:98]
  wire [63:0] _aluWbData_T_6 = 2'h2 == exInsts_0_src_b ? csr_io_common_io_out : alu_io_r; // @[Mux.scala 80:57]
  wire [63:0] aluWbData = exInsts_0_write_src == 2'h3 | exInsts_0_next_pc != 4'h0 ? {{32'd0}, _exReBranchPC_T_3} :
    _aluWbData_T_6; // @[Backend.scala 423:19]
  wire [63:0] _GEN_24 = exInsts_0_rd == issueInsts_0_rs1 ? aluWbData : _GEN_20; // @[Backend.scala 197:49 Backend.scala 198:22]
  wire [63:0] _GEN_25 = exInsts_0_rd == issueInsts_0_rs2 ? aluWbData : _GEN_21; // @[Backend.scala 200:49 Backend.scala 201:22]
  wire [63:0] _GEN_26 = exInsts_0_rd == issueInsts_1_rs1 ? aluWbData : _GEN_22; // @[Backend.scala 197:49 Backend.scala 198:22]
  wire [63:0] _GEN_27 = exInsts_0_rd == issueInsts_1_rs2 ? aluWbData : _GEN_23; // @[Backend.scala 200:49 Backend.scala 201:22]
  wire [63:0] _GEN_28 = exInstsValid_0 & exInsts_0_write_dest & exInsts_0_rd != 5'h0 ? _GEN_24 : _GEN_20; // @[Backend.scala 195:96]
  wire [63:0] _GEN_29 = exInstsValid_0 & exInsts_0_write_dest & exInsts_0_rd != 5'h0 ? _GEN_25 : _GEN_21; // @[Backend.scala 195:96]
  wire [63:0] _GEN_30 = exInstsValid_0 & exInsts_0_write_dest & exInsts_0_rd != 5'h0 ? _GEN_26 : _GEN_22; // @[Backend.scala 195:96]
  wire [63:0] _GEN_31 = exInstsValid_0 & exInsts_0_write_dest & exInsts_0_rd != 5'h0 ? _GEN_27 : _GEN_23; // @[Backend.scala 195:96]
  wire [63:0] _GEN_32 = exInsts_1_rd == issueInsts_0_rs1 ? mdu_io_resp_r : _GEN_28; // @[Backend.scala 207:49 Backend.scala 208:22]
  wire [63:0] _GEN_33 = exInsts_1_rd == issueInsts_0_rs2 ? mdu_io_resp_r : _GEN_29; // @[Backend.scala 210:49 Backend.scala 211:22]
  wire [63:0] _GEN_34 = exInsts_1_rd == issueInsts_1_rs1 ? mdu_io_resp_r : _GEN_30; // @[Backend.scala 207:49 Backend.scala 208:22]
  wire [63:0] _GEN_35 = exInsts_1_rd == issueInsts_1_rs2 ? mdu_io_resp_r : _GEN_31; // @[Backend.scala 210:49 Backend.scala 211:22]
  wire [31:0] genImm_1_hi_hi = exInsts_1_imm[19] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_1_T_5 = {genImm_1_hi_hi,exInsts_1_imm,12'h0}; // @[Cat.scala 30:58]
  wire [43:0] genImm_1_hi_1 = exInsts_1_imm[19] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _genImm_1_T_8 = {genImm_1_hi_1,exInsts_1_imm}; // @[Cat.scala 30:58]
  wire [63:0] genImm_1 = exInsts_1_alu_op == 5'ha | exInsts_1_src_a == 2'h2 ? _genImm_1_T_5 : _genImm_1_T_8; // @[Backend.scala 54:8]
  wire [2:0] _exInstsValid_0_T = {issueArbiter_io_issue_fu_valid_2,issueArbiter_io_issue_fu_valid_1,
    issueArbiter_io_issue_fu_valid_0}; // @[Backend.scala 254:57]
  wire  nop_ysyx_print = 1'h0; // @[Backend.scala 26:19 Backend.scala 47:22]
  wire [31:0] issueInsts_0_pc = issueQueue_io_dout_0_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  wire [63:0] issueRss_0 = issueArbiter_io_rss_out_0; // @[Backend.scala 66:26 Backend.scala 172:31]
  wire [63:0] issueRts_0 = issueArbiter_io_rts_out_0; // @[Backend.scala 67:26 Backend.scala 173:31]
  wire [63:0] issueRss_1 = issueArbiter_io_rss_out_1; // @[Backend.scala 66:26 Backend.scala 172:31]
  wire [63:0] issueRts_1 = issueArbiter_io_rts_out_1; // @[Backend.scala 67:26 Backend.scala 173:31]
  wire [63:0] issueRss_2 = issueArbiter_io_rss_out_2; // @[Backend.scala 66:26 Backend.scala 172:31]
  wire [63:0] issueRts_2 = issueArbiter_io_rts_out_2; // @[Backend.scala 67:26 Backend.scala 173:31]
  wire  mduValid = exInstsValid_1 & _aluValid_T; // @[Backend.scala 280:33]
  wire [63:0] _alu_io_a_T = {59'h0,exInsts_0_rs1}; // @[Cat.scala 30:58]
  wire [63:0] _alu_io_a_T_2 = 2'h2 == exInsts_0_src_a ? {{32'd0}, exInsts_0_pc} : exFwdRsData_0; // @[Mux.scala 80:57]
  wire  ldMisaligned = exInsts_2_write_dest & memMisaligned; // @[Backend.scala 309:62]
  wire  stMisaligned = ~exInsts_2_write_dest & memMisaligned; // @[Backend.scala 310:62]
  wire [1:0] _exMemReq_memReq_mtype_T_1 = 3'h1 == exInsts_2_mem_width ? 2'h0 : 2'h2; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_3 = 3'h0 == exInsts_2_mem_width ? 2'h0 : _exMemReq_memReq_mtype_T_1; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_5 = 3'h2 == exInsts_2_mem_width ? 2'h1 : _exMemReq_memReq_mtype_T_3; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_7 = 3'h3 == exInsts_2_mem_width ? 2'h1 : _exMemReq_memReq_mtype_T_5; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_9 = 3'h4 == exInsts_2_mem_width ? 2'h2 : _exMemReq_memReq_mtype_T_7; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_11 = 3'h5 == exInsts_2_mem_width ? 2'h3 : _exMemReq_memReq_mtype_T_9; // @[Mux.scala 80:57]
  wire [1:0] _exMemReq_memReq_mtype_T_13 = 3'h6 == exInsts_2_mem_width ? 2'h2 : _exMemReq_memReq_mtype_T_11; // @[Mux.scala 80:57]
  wire [31:0] exMemReq_addr = ldstAddr[31:0]; // @[Backend.scala 339:22 Backend.scala 344:18]
  wire  _GEN_218 = isExPCJump ? _bpuErrpr_T_7 | ~exInsts_0_predict_taken | |jumpPc[1:0] : exCsrValid; // @[Backend.scala 393:29 Backend.scala 394:16]
  wire  _GEN_220 = isExPCBr ? reBranchBrTaken ^ exInsts_0_predict_taken | reBranchBrTaken & (_bpuErrpr_T_2 | |brPC[1:0])
     : _GEN_218; // @[Backend.scala 370:21 Backend.scala 381:16]
  wire  reBranch = exInstsTrueValid_0 & _GEN_220; // @[Backend.scala 369:29 Backend.scala 362:12]
  wire  exInstsTrueValid_1 = mduValid & ~mduExptMask; // @[Backend.scala 415:35]
  wire  _GEN_230 = _issueQueue_io_deqReq_T & bpuV; // @[Backend.scala 462:26 Backend.scala 464:12 Backend.scala 485:12]
  wire [63:0] _GEN_306 = _issueQueue_io_deqReq_T ? exReBranchPC : {{32'd0}, reBranchPC}; // @[Backend.scala 462:26 Backend.scala 480:16 Backend.scala 124:29]
  wire [63:0] _GEN_386 = io_fb_bmfs_redirect_kill ? {{32'd0}, reBranchPC} : _GEN_306; // @[Backend.scala 455:17 Backend.scala 124:29]
  wire [63:0] _io_fb_bmfs_redirect_pc_T = csr_io_event_io_except_kill ? csr_io_event_io_redirect_pc : {{32'd0},
    reBranchPC}; // @[Backend.scala 489:34]
  wire  wbExcepts_0 = |wbInsts__0_pc[1:0]; // @[Backend.scala 522:39]
  wire  _regFile_io_wen_vec_0_T_1 = ~wbExcepts_0; // @[Backend.scala 498:68]
  wire  _regFile_io_wen_vec_0_T_2 = wbInsts__0_write_dest & ~wbExcepts_0; // @[Backend.scala 498:65]
  wire  wbExcepts_1 = |wbInsts__1_pc[1:0]; // @[Backend.scala 523:39]
  wire  _regFile_io_wen_vec_0_T_5 = ~wbExcepts_1; // @[Backend.scala 499:70]
  wire  _regFile_io_wen_vec_0_T_6 = _T_9 & ~wbExcepts_1; // @[Backend.scala 499:67]
  wire  wbLdMaReal = wbInstsValid_2 & wbLdMa; // @[Backend.scala 515:39]
  wire  _regFile_io_wen_vec_1_T_1 = ~wbLdMaReal; // @[Backend.scala 505:68]
  wire  _regFile_io_wen_vec_1_T_2 = wbInsts__2_write_dest & ~wbLdMaReal; // @[Backend.scala 505:65]
  wire  csrWbValid = wbInsts__0_next_pc == 4'h0 & wbInsts__0_alu_mdu_lsu == 2'h0; // @[Backend.scala 513:62]
  wire  wbALUSysReal = wbInsts__0_next_pc == 4'h5 & wbInstsValid_0; // @[Backend.scala 517:63]
  wire  wbALUBpReal = wbInsts__0_next_pc == 4'h8 & wbInstsValid_0; // @[Backend.scala 518:64]
  wire  illegal = wbInsts__0_illegal & wbInstsValid_0; // @[Backend.scala 519:42]
  wire  wbFetchMaReal = wbExcepts_0 & wbInstsValid_0; // @[Backend.scala 520:47]
  wire [2:0] _wb_deal_with_int_T = {wbInstsValid_2,wbInstsValid_1,wbInstsValid_0}; // @[Backend.scala 542:61]
  wire  wb_deal_with_int = wbInterruptd & |_wb_deal_with_int_T & exInterruptd; // @[Backend.scala 542:91]
  wire [63:0] wb_pc_0 = wbInstsValid_0 ? {{32'd0}, wbInsts__0_pc} : 64'hffffffffffffffff; // @[Backend.scala 545:20]
  wire [63:0] wb_pc_1 = wbInstsValid_1 ? {{32'd0}, wbInsts__1_pc} : 64'hffffffffffffffff; // @[Backend.scala 545:20]
  wire [63:0] wb_pc_2 = wbInstsValid_2 ? {{32'd0}, wbInsts__2_pc} : 64'hffffffffffffffff; // @[Backend.scala 545:20]
  wire [63:0] _wb_pc_min_T_2 = wb_pc_0 < wb_pc_2 ? wb_pc_0 : wb_pc_2; // @[Backend.scala 547:8]
  wire [63:0] _wb_pc_min_T_4 = wb_pc_1 < wb_pc_2 ? wb_pc_1 : wb_pc_2; // @[Backend.scala 548:8]
  wire [63:0] wb_pc_min = wb_pc_0 < wb_pc_1 ? _wb_pc_min_T_2 : _wb_pc_min_T_4; // @[Backend.scala 546:22]
  wire [31:0] _csr_io_event_io_epc_T_2 = wbALUSysReal | wbALUBpReal | illegal ? wbInsts__0_pc : wbInsts__1_pc; // @[Backend.scala 566:8]
  wire [31:0] _csr_io_event_io_bad_address_T = wbFetchMaReal ? wbInsts__0_pc : wbMisalignedAddr; // @[Backend.scala 567:37]
  reg [31:0] bufInsts0_pc; // @[Backend.scala 590:59]
  reg [31:0] bufInsts0_inst; // @[Backend.scala 590:59]
  reg  bufInstsValid0; // @[Backend.scala 590:74]
  reg [1:0] bufInstsOrder0; // @[Backend.scala 590:87]
  reg  REG; // @[Backend.scala 591:33]
  reg  tmp_REG; // @[Backend.scala 598:28]
  reg  REG_1; // @[Backend.scala 599:26]
  wire  _tmp_T_13 = wbInstsValid_1 & _issueQueue_io_deqReq_T; // @[Backend.scala 598:112]
  wire  _tmp_T_14 = |wbInsts__1_inst; // @[Backend.scala 598:147]
  reg  REG_2; // @[Backend.scala 600:19]
  wire  _tmp_T_21 = wbInstsValid_2 & _issueQueue_io_deqReq_T; // @[Backend.scala 598:112]
  wire  _tmp_T_22 = |wbInsts__2_inst; // @[Backend.scala 598:147]
  reg  REG_3; // @[Backend.scala 600:19]
  reg  tmp_REG_3; // @[Backend.scala 603:28]
  reg [31:0] REG_4; // @[Backend.scala 604:26]
  reg [31:0] REG_5; // @[Backend.scala 605:19]
  reg [31:0] REG_6; // @[Backend.scala 605:19]
  reg  tmp_REG_6; // @[Backend.scala 608:28]
  reg [1:0] REG_7; // @[Backend.scala 609:26]
  reg [1:0] REG_8; // @[Backend.scala 610:19]
  reg [1:0] REG_9; // @[Backend.scala 610:19]
  reg  tmp_REG_9; // @[Backend.scala 613:28]
  reg [31:0] REG_10; // @[Backend.scala 614:26]
  reg [31:0] REG_11; // @[Backend.scala 615:19]
  reg [31:0] REG_12; // @[Backend.scala 615:19]
  reg  REG_13; // @[Backend.scala 617:72]
  reg  REG_14; // @[Backend.scala 623:60]
  reg  REG_15; // @[Backend.scala 623:60]
  reg  REG_16; // @[Backend.scala 623:60]
  reg [63:0] instret; // @[Backend.scala 627:26]
  reg [63:0] counter; // @[Backend.scala 628:26]
  reg [63:0] dstall; // @[Backend.scala 629:25]
  reg [63:0] istall; // @[Backend.scala 631:25]
  reg [63:0] mduStall; // @[Backend.scala 632:27]
  reg [63:0] common; // @[Backend.scala 633:25]
  wire [63:0] _GEN_412 = {{63'd0}, dcacheStall}; // @[Backend.scala 635:22]
  wire [63:0] _dstall_T_2 = dstall + _GEN_412; // @[Backend.scala 635:22]
  wire [63:0] _GEN_413 = {{63'd0}, icache_stall}; // @[Backend.scala 636:22]
  wire [63:0] _istall_T_2 = istall + _GEN_413; // @[Backend.scala 636:22]
  wire  _common_T = dcacheStall & icache_stall; // @[Backend.scala 637:40]
  wire [63:0] _GEN_414 = {{63'd0}, _common_T}; // @[Backend.scala 637:22]
  wire [63:0] _common_T_3 = common + _GEN_414; // @[Backend.scala 637:22]
  wire [63:0] _counter_T_1 = counter + 64'h1; // @[Backend.scala 638:24]
  wire  _instret_T_1 = wbInstsValid_0 & _regFile_io_wen_vec_0_T_1; // @[Backend.scala 639:66]
  wire [63:0] _GEN_415 = {{63'd0}, _instret_T_1}; // @[Backend.scala 639:47]
  wire [63:0] _instret_T_3 = instret + _GEN_415; // @[Backend.scala 639:47]
  wire  _instret_T_5 = wbInstsValid_1 & _regFile_io_wen_vec_0_T_5; // @[Backend.scala 639:110]
  wire [63:0] _GEN_416 = {{63'd0}, _instret_T_5}; // @[Backend.scala 639:91]
  wire [63:0] _instret_T_7 = _instret_T_3 + _GEN_416; // @[Backend.scala 639:91]
  wire  _instret_T_9 = wbInstsValid_2 & _regFile_io_wen_vec_1_T_1; // @[Backend.scala 639:154]
  wire [63:0] _GEN_417 = {{63'd0}, _instret_T_9}; // @[Backend.scala 639:135]
  wire [63:0] _instret_T_11 = _instret_T_7 + _GEN_417; // @[Backend.scala 639:135]
  wire [63:0] _GEN_418 = {{63'd0}, _stall_i_T}; // @[Backend.scala 640:26]
  wire [63:0] _mduStall_T_2 = mduStall + _GEN_418; // @[Backend.scala 640:26]
  wire  _WIRE__0 = REG_1; // @[Backend.scala 597:34 Backend.scala 597:34]
  wire  _WIRE__1 = REG_2; // @[Backend.scala 597:34 Backend.scala 597:34]
  wire  _WIRE__2 = REG_3; // @[Backend.scala 597:34 Backend.scala 597:34]
  wire [31:0] _WIRE_1_0 = REG_4; // @[Backend.scala 602:34 Backend.scala 602:34]
  wire [31:0] _WIRE_1_1 = REG_5; // @[Backend.scala 602:34 Backend.scala 602:34]
  wire [31:0] _WIRE_1_2 = REG_6; // @[Backend.scala 602:34 Backend.scala 602:34]
  wire [1:0] _WIRE_2_0 = REG_7; // @[Backend.scala 607:34 Backend.scala 607:34]
  wire [1:0] _WIRE_2_1 = REG_8; // @[Backend.scala 607:34 Backend.scala 607:34]
  wire [1:0] _WIRE_2_2 = REG_9; // @[Backend.scala 607:34 Backend.scala 607:34]
  wire [31:0] _WIRE_3_0 = REG_10; // @[Backend.scala 612:34 Backend.scala 612:34]
  wire [31:0] _WIRE_3_1 = REG_11; // @[Backend.scala 612:34 Backend.scala 612:34]
  wire [31:0] _WIRE_3_2 = REG_12; // @[Backend.scala 612:34 Backend.scala 612:34]
  wire  _WIRE_4_0 = 1'h0; // @[Backend.scala 617:34 Backend.scala 617:34]
  wire  _WIRE_4_1 = 1'h0; // @[Backend.scala 617:34 Backend.scala 617:34]
  wire  _WIRE_4_2 = REG_13; // @[Backend.scala 617:34 Backend.scala 617:34]
  wire  _WIRE_5_0 = REG_14; // @[Backend.scala 623:34 Backend.scala 623:34]
  wire  _WIRE_5_1 = REG_15; // @[Backend.scala 623:34 Backend.scala 623:34]
  wire  _WIRE_5_2 = REG_16; // @[Backend.scala 623:34 Backend.scala 623:34]
  ALU alu ( // @[Backend.scala 59:28]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_aluOp(alu_io_aluOp),
    .io_aluExpand(alu_io_aluExpand),
    .io_aluCsr(alu_io_aluCsr),
    .io_csr(alu_io_csr),
    .io_r(alu_io_r),
    .io_zero(alu_io_zero)
  );
  MDU mdu ( // @[Backend.scala 60:28]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_kill(mdu_io_kill),
    .io_req_valid(mdu_io_req_valid),
    .io_req_op(mdu_io_req_op),
    .io_req_expand(mdu_io_req_expand),
    .io_req_in1(mdu_io_req_in1),
    .io_req_in2(mdu_io_req_in2),
    .io_resp_r(mdu_io_resp_r),
    .io_resp_valid(mdu_io_resp_valid)
  );
  FIFO issueQueue ( // @[Backend.scala 68:28]
    .clock(issueQueue_clock),
    .reset(issueQueue_reset),
    .io_dout_0_illegal(issueQueue_io_dout_0_illegal),
    .io_dout_0_next_pc(issueQueue_io_dout_0_next_pc),
    .io_dout_0_alu_mdu_lsu(issueQueue_io_dout_0_alu_mdu_lsu),
    .io_dout_0_branch_type(issueQueue_io_dout_0_branch_type),
    .io_dout_0_src_a(issueQueue_io_dout_0_src_a),
    .io_dout_0_src_b(issueQueue_io_dout_0_src_b),
    .io_dout_0_write_dest(issueQueue_io_dout_0_write_dest),
    .io_dout_0_alu_op(issueQueue_io_dout_0_alu_op),
    .io_dout_0_alu_expand(issueQueue_io_dout_0_alu_expand),
    .io_dout_0_mem_width(issueQueue_io_dout_0_mem_width),
    .io_dout_0_write_src(issueQueue_io_dout_0_write_src),
    .io_dout_0_rs1(issueQueue_io_dout_0_rs1),
    .io_dout_0_rs2(issueQueue_io_dout_0_rs2),
    .io_dout_0_rd(issueQueue_io_dout_0_rd),
    .io_dout_0_imm(issueQueue_io_dout_0_imm),
    .io_dout_0_pc(issueQueue_io_dout_0_pc),
    .io_dout_0_predict_taken(issueQueue_io_dout_0_predict_taken),
    .io_dout_0_target_pc(issueQueue_io_dout_0_target_pc),
    .io_dout_0_ysyx_debug(issueQueue_io_dout_0_ysyx_debug),
    .io_dout_0_ysyx_print(issueQueue_io_dout_0_ysyx_print),
    .io_dout_0_inst(issueQueue_io_dout_0_inst),
    .io_dout_1_illegal(issueQueue_io_dout_1_illegal),
    .io_dout_1_next_pc(issueQueue_io_dout_1_next_pc),
    .io_dout_1_alu_mdu_lsu(issueQueue_io_dout_1_alu_mdu_lsu),
    .io_dout_1_branch_type(issueQueue_io_dout_1_branch_type),
    .io_dout_1_src_a(issueQueue_io_dout_1_src_a),
    .io_dout_1_src_b(issueQueue_io_dout_1_src_b),
    .io_dout_1_write_dest(issueQueue_io_dout_1_write_dest),
    .io_dout_1_alu_op(issueQueue_io_dout_1_alu_op),
    .io_dout_1_alu_expand(issueQueue_io_dout_1_alu_expand),
    .io_dout_1_mem_width(issueQueue_io_dout_1_mem_width),
    .io_dout_1_write_src(issueQueue_io_dout_1_write_src),
    .io_dout_1_rs1(issueQueue_io_dout_1_rs1),
    .io_dout_1_rs2(issueQueue_io_dout_1_rs2),
    .io_dout_1_rd(issueQueue_io_dout_1_rd),
    .io_dout_1_imm(issueQueue_io_dout_1_imm),
    .io_dout_1_pc(issueQueue_io_dout_1_pc),
    .io_dout_1_predict_taken(issueQueue_io_dout_1_predict_taken),
    .io_dout_1_target_pc(issueQueue_io_dout_1_target_pc),
    .io_dout_1_ysyx_debug(issueQueue_io_dout_1_ysyx_debug),
    .io_dout_1_ysyx_print(issueQueue_io_dout_1_ysyx_print),
    .io_dout_1_inst(issueQueue_io_dout_1_inst),
    .io_enqStep(issueQueue_io_enqStep),
    .io_enqReq(issueQueue_io_enqReq),
    .io_deqStep(issueQueue_io_deqStep),
    .io_deqReq(issueQueue_io_deqReq),
    .io_din_0_illegal(issueQueue_io_din_0_illegal),
    .io_din_0_next_pc(issueQueue_io_din_0_next_pc),
    .io_din_0_alu_mdu_lsu(issueQueue_io_din_0_alu_mdu_lsu),
    .io_din_0_branch_type(issueQueue_io_din_0_branch_type),
    .io_din_0_src_a(issueQueue_io_din_0_src_a),
    .io_din_0_src_b(issueQueue_io_din_0_src_b),
    .io_din_0_write_dest(issueQueue_io_din_0_write_dest),
    .io_din_0_alu_op(issueQueue_io_din_0_alu_op),
    .io_din_0_alu_expand(issueQueue_io_din_0_alu_expand),
    .io_din_0_mem_width(issueQueue_io_din_0_mem_width),
    .io_din_0_write_src(issueQueue_io_din_0_write_src),
    .io_din_0_rs1(issueQueue_io_din_0_rs1),
    .io_din_0_rs2(issueQueue_io_din_0_rs2),
    .io_din_0_rd(issueQueue_io_din_0_rd),
    .io_din_0_imm(issueQueue_io_din_0_imm),
    .io_din_0_pc(issueQueue_io_din_0_pc),
    .io_din_0_predict_taken(issueQueue_io_din_0_predict_taken),
    .io_din_0_target_pc(issueQueue_io_din_0_target_pc),
    .io_din_0_ysyx_debug(issueQueue_io_din_0_ysyx_debug),
    .io_din_0_ysyx_print(issueQueue_io_din_0_ysyx_print),
    .io_din_0_inst(issueQueue_io_din_0_inst),
    .io_din_1_illegal(issueQueue_io_din_1_illegal),
    .io_din_1_next_pc(issueQueue_io_din_1_next_pc),
    .io_din_1_alu_mdu_lsu(issueQueue_io_din_1_alu_mdu_lsu),
    .io_din_1_branch_type(issueQueue_io_din_1_branch_type),
    .io_din_1_src_a(issueQueue_io_din_1_src_a),
    .io_din_1_src_b(issueQueue_io_din_1_src_b),
    .io_din_1_write_dest(issueQueue_io_din_1_write_dest),
    .io_din_1_alu_op(issueQueue_io_din_1_alu_op),
    .io_din_1_alu_expand(issueQueue_io_din_1_alu_expand),
    .io_din_1_mem_width(issueQueue_io_din_1_mem_width),
    .io_din_1_write_src(issueQueue_io_din_1_write_src),
    .io_din_1_rs1(issueQueue_io_din_1_rs1),
    .io_din_1_rs2(issueQueue_io_din_1_rs2),
    .io_din_1_rd(issueQueue_io_din_1_rd),
    .io_din_1_imm(issueQueue_io_din_1_imm),
    .io_din_1_pc(issueQueue_io_din_1_pc),
    .io_din_1_predict_taken(issueQueue_io_din_1_predict_taken),
    .io_din_1_target_pc(issueQueue_io_din_1_target_pc),
    .io_din_1_ysyx_debug(issueQueue_io_din_1_ysyx_debug),
    .io_din_1_ysyx_print(issueQueue_io_din_1_ysyx_print),
    .io_din_1_inst(issueQueue_io_din_1_inst),
    .io_flush(issueQueue_io_flush),
    .io_sufficient(issueQueue_io_sufficient),
    .io_items(issueQueue_io_items)
  );
  IssueArbiter issueArbiter ( // @[Backend.scala 69:28]
    .io_insts_in_0_illegal(issueArbiter_io_insts_in_0_illegal),
    .io_insts_in_0_next_pc(issueArbiter_io_insts_in_0_next_pc),
    .io_insts_in_0_alu_mdu_lsu(issueArbiter_io_insts_in_0_alu_mdu_lsu),
    .io_insts_in_0_branch_type(issueArbiter_io_insts_in_0_branch_type),
    .io_insts_in_0_src_a(issueArbiter_io_insts_in_0_src_a),
    .io_insts_in_0_src_b(issueArbiter_io_insts_in_0_src_b),
    .io_insts_in_0_write_dest(issueArbiter_io_insts_in_0_write_dest),
    .io_insts_in_0_alu_op(issueArbiter_io_insts_in_0_alu_op),
    .io_insts_in_0_alu_expand(issueArbiter_io_insts_in_0_alu_expand),
    .io_insts_in_0_mem_width(issueArbiter_io_insts_in_0_mem_width),
    .io_insts_in_0_write_src(issueArbiter_io_insts_in_0_write_src),
    .io_insts_in_0_rs1(issueArbiter_io_insts_in_0_rs1),
    .io_insts_in_0_rs2(issueArbiter_io_insts_in_0_rs2),
    .io_insts_in_0_rd(issueArbiter_io_insts_in_0_rd),
    .io_insts_in_0_imm(issueArbiter_io_insts_in_0_imm),
    .io_insts_in_0_pc(issueArbiter_io_insts_in_0_pc),
    .io_insts_in_0_predict_taken(issueArbiter_io_insts_in_0_predict_taken),
    .io_insts_in_0_target_pc(issueArbiter_io_insts_in_0_target_pc),
    .io_insts_in_0_ysyx_debug(issueArbiter_io_insts_in_0_ysyx_debug),
    .io_insts_in_0_ysyx_print(issueArbiter_io_insts_in_0_ysyx_print),
    .io_insts_in_0_inst(issueArbiter_io_insts_in_0_inst),
    .io_insts_in_1_illegal(issueArbiter_io_insts_in_1_illegal),
    .io_insts_in_1_next_pc(issueArbiter_io_insts_in_1_next_pc),
    .io_insts_in_1_alu_mdu_lsu(issueArbiter_io_insts_in_1_alu_mdu_lsu),
    .io_insts_in_1_branch_type(issueArbiter_io_insts_in_1_branch_type),
    .io_insts_in_1_src_a(issueArbiter_io_insts_in_1_src_a),
    .io_insts_in_1_src_b(issueArbiter_io_insts_in_1_src_b),
    .io_insts_in_1_write_dest(issueArbiter_io_insts_in_1_write_dest),
    .io_insts_in_1_alu_op(issueArbiter_io_insts_in_1_alu_op),
    .io_insts_in_1_alu_expand(issueArbiter_io_insts_in_1_alu_expand),
    .io_insts_in_1_mem_width(issueArbiter_io_insts_in_1_mem_width),
    .io_insts_in_1_write_src(issueArbiter_io_insts_in_1_write_src),
    .io_insts_in_1_rs1(issueArbiter_io_insts_in_1_rs1),
    .io_insts_in_1_rs2(issueArbiter_io_insts_in_1_rs2),
    .io_insts_in_1_rd(issueArbiter_io_insts_in_1_rd),
    .io_insts_in_1_imm(issueArbiter_io_insts_in_1_imm),
    .io_insts_in_1_pc(issueArbiter_io_insts_in_1_pc),
    .io_insts_in_1_predict_taken(issueArbiter_io_insts_in_1_predict_taken),
    .io_insts_in_1_target_pc(issueArbiter_io_insts_in_1_target_pc),
    .io_insts_in_1_ysyx_debug(issueArbiter_io_insts_in_1_ysyx_debug),
    .io_insts_in_1_ysyx_print(issueArbiter_io_insts_in_1_ysyx_print),
    .io_insts_in_1_inst(issueArbiter_io_insts_in_1_inst),
    .io_queue_items(issueArbiter_io_queue_items),
    .io_ld_dest_ex(issueArbiter_io_ld_dest_ex),
    .io_rss_in_0(issueArbiter_io_rss_in_0),
    .io_rss_in_1(issueArbiter_io_rss_in_1),
    .io_rts_in_0(issueArbiter_io_rts_in_0),
    .io_rts_in_1(issueArbiter_io_rts_in_1),
    .io_rss_out_0(issueArbiter_io_rss_out_0),
    .io_rss_out_1(issueArbiter_io_rss_out_1),
    .io_rss_out_2(issueArbiter_io_rss_out_2),
    .io_rts_out_0(issueArbiter_io_rts_out_0),
    .io_rts_out_1(issueArbiter_io_rts_out_1),
    .io_rts_out_2(issueArbiter_io_rts_out_2),
    .io_insts_out_0_illegal(issueArbiter_io_insts_out_0_illegal),
    .io_insts_out_0_next_pc(issueArbiter_io_insts_out_0_next_pc),
    .io_insts_out_0_alu_mdu_lsu(issueArbiter_io_insts_out_0_alu_mdu_lsu),
    .io_insts_out_0_branch_type(issueArbiter_io_insts_out_0_branch_type),
    .io_insts_out_0_src_a(issueArbiter_io_insts_out_0_src_a),
    .io_insts_out_0_src_b(issueArbiter_io_insts_out_0_src_b),
    .io_insts_out_0_write_dest(issueArbiter_io_insts_out_0_write_dest),
    .io_insts_out_0_alu_op(issueArbiter_io_insts_out_0_alu_op),
    .io_insts_out_0_alu_expand(issueArbiter_io_insts_out_0_alu_expand),
    .io_insts_out_0_write_src(issueArbiter_io_insts_out_0_write_src),
    .io_insts_out_0_rs1(issueArbiter_io_insts_out_0_rs1),
    .io_insts_out_0_rd(issueArbiter_io_insts_out_0_rd),
    .io_insts_out_0_imm(issueArbiter_io_insts_out_0_imm),
    .io_insts_out_0_pc(issueArbiter_io_insts_out_0_pc),
    .io_insts_out_0_predict_taken(issueArbiter_io_insts_out_0_predict_taken),
    .io_insts_out_0_target_pc(issueArbiter_io_insts_out_0_target_pc),
    .io_insts_out_0_ysyx_debug(issueArbiter_io_insts_out_0_ysyx_debug),
    .io_insts_out_0_ysyx_print(issueArbiter_io_insts_out_0_ysyx_print),
    .io_insts_out_0_inst(issueArbiter_io_insts_out_0_inst),
    .io_insts_out_1_src_a(issueArbiter_io_insts_out_1_src_a),
    .io_insts_out_1_src_b(issueArbiter_io_insts_out_1_src_b),
    .io_insts_out_1_write_dest(issueArbiter_io_insts_out_1_write_dest),
    .io_insts_out_1_alu_op(issueArbiter_io_insts_out_1_alu_op),
    .io_insts_out_1_alu_expand(issueArbiter_io_insts_out_1_alu_expand),
    .io_insts_out_1_rd(issueArbiter_io_insts_out_1_rd),
    .io_insts_out_1_imm(issueArbiter_io_insts_out_1_imm),
    .io_insts_out_1_pc(issueArbiter_io_insts_out_1_pc),
    .io_insts_out_1_ysyx_print(issueArbiter_io_insts_out_1_ysyx_print),
    .io_insts_out_1_inst(issueArbiter_io_insts_out_1_inst),
    .io_insts_out_2_src_a(issueArbiter_io_insts_out_2_src_a),
    .io_insts_out_2_write_dest(issueArbiter_io_insts_out_2_write_dest),
    .io_insts_out_2_alu_op(issueArbiter_io_insts_out_2_alu_op),
    .io_insts_out_2_mem_width(issueArbiter_io_insts_out_2_mem_width),
    .io_insts_out_2_rd(issueArbiter_io_insts_out_2_rd),
    .io_insts_out_2_imm(issueArbiter_io_insts_out_2_imm),
    .io_insts_out_2_pc(issueArbiter_io_insts_out_2_pc),
    .io_insts_out_2_ysyx_print(issueArbiter_io_insts_out_2_ysyx_print),
    .io_insts_out_2_inst(issueArbiter_io_insts_out_2_inst),
    .io_issue_num(issueArbiter_io_issue_num),
    .io_issue_fu_valid_0(issueArbiter_io_issue_fu_valid_0),
    .io_issue_fu_valid_1(issueArbiter_io_issue_fu_valid_1),
    .io_issue_fu_valid_2(issueArbiter_io_issue_fu_valid_2),
    .io_insts_order_0(issueArbiter_io_insts_order_0),
    .io_insts_order_1(issueArbiter_io_insts_order_1),
    .io_insts_order_2(issueArbiter_io_insts_order_2)
  );
  RegFile regFile ( // @[Backend.scala 131:32]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_rs_addr_vec_0(regFile_io_rs_addr_vec_0),
    .io_rs_addr_vec_1(regFile_io_rs_addr_vec_1),
    .io_rs_addr_vec_2(regFile_io_rs_addr_vec_2),
    .io_rs_addr_vec_3(regFile_io_rs_addr_vec_3),
    .io_rs_data_vec_0(regFile_io_rs_data_vec_0),
    .io_rs_data_vec_1(regFile_io_rs_data_vec_1),
    .io_rs_data_vec_2(regFile_io_rs_data_vec_2),
    .io_rs_data_vec_3(regFile_io_rs_data_vec_3),
    .io_wen_vec_0(regFile_io_wen_vec_0),
    .io_wen_vec_1(regFile_io_wen_vec_1),
    .io_rd_addr_vec_0(regFile_io_rd_addr_vec_0),
    .io_rd_addr_vec_1(regFile_io_rd_addr_vec_1),
    .io_rd_data_vec_0(regFile_io_rd_data_vec_0),
    .io_rd_data_vec_1(regFile_io_rd_data_vec_1),
    .difftestSaddr(regFile_difftestSaddr),
    ._WIRE_0_0(regFile__WIRE_0_0),
    ._WIRE_0_1(regFile__WIRE_0_1),
    ._WIRE_0_2(regFile__WIRE_0_2),
    ._WIRE_0_3(regFile__WIRE_0_3),
    ._WIRE_0_4(regFile__WIRE_0_4),
    ._WIRE_0_5(regFile__WIRE_0_5),
    ._WIRE_0_6(regFile__WIRE_0_6),
    ._WIRE_0_7(regFile__WIRE_0_7),
    ._WIRE_0_8(regFile__WIRE_0_8),
    ._WIRE_0_9(regFile__WIRE_0_9),
    ._WIRE_0_10(regFile__WIRE_0_10),
    ._WIRE_0_11(regFile__WIRE_0_11),
    ._WIRE_0_12(regFile__WIRE_0_12),
    ._WIRE_0_13(regFile__WIRE_0_13),
    ._WIRE_0_14(regFile__WIRE_0_14),
    ._WIRE_0_15(regFile__WIRE_0_15),
    ._WIRE_0_16(regFile__WIRE_0_16),
    ._WIRE_0_17(regFile__WIRE_0_17),
    ._WIRE_0_18(regFile__WIRE_0_18),
    ._WIRE_0_19(regFile__WIRE_0_19),
    ._WIRE_0_20(regFile__WIRE_0_20),
    ._WIRE_0_21(regFile__WIRE_0_21),
    ._WIRE_0_22(regFile__WIRE_0_22),
    ._WIRE_0_23(regFile__WIRE_0_23),
    ._WIRE_0_24(regFile__WIRE_0_24),
    ._WIRE_0_25(regFile__WIRE_0_25),
    ._WIRE_0_26(regFile__WIRE_0_26),
    ._WIRE_0_27(regFile__WIRE_0_27),
    ._WIRE_0_28(regFile__WIRE_0_28),
    ._WIRE_0_29(regFile__WIRE_0_29),
    ._WIRE_0_30(regFile__WIRE_0_30),
    ._WIRE_0_31(regFile__WIRE_0_31),
    .difftestSval(regFile_difftestSval),
    .difftestSync(regFile_difftestSync)
  );
  CSR csr ( // @[Backend.scala 132:32]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_common_io_in(csr_io_common_io_in),
    .io_common_io_wen(csr_io_common_io_wen),
    .io_common_io_num(csr_io_common_io_num),
    .io_common_io_out(csr_io_common_io_out),
    .io_event_io_exception_vec_2(csr_io_event_io_exception_vec_2),
    .io_event_io_exception_vec_3(csr_io_event_io_exception_vec_3),
    .io_event_io_exception_vec_4(csr_io_event_io_exception_vec_4),
    .io_event_io_exception_vec_6(csr_io_event_io_exception_vec_6),
    .io_event_io_deal_with_int(csr_io_event_io_deal_with_int),
    .io_event_io_is_mret(csr_io_event_io_is_mret),
    .io_event_io_is_sret(csr_io_event_io_is_sret),
    .io_event_io_is_ecall(csr_io_event_io_is_ecall),
    .io_event_io_bad_address(csr_io_event_io_bad_address),
    .io_event_io_epc(csr_io_event_io_epc),
    .io_event_io_call_for_int(csr_io_event_io_call_for_int),
    .io_event_io_except_kill(csr_io_event_io_except_kill),
    .io_event_io_redirect_pc(csr_io_event_io_redirect_pc),
    .csrs_0_mstatus(csr_csrs_0_mstatus),
    .csrs_0_sstatus(csr_csrs_0_sstatus),
    .csrs_0_mepc(csr_csrs_0_mepc),
    .csrs_0_sepc(csr_csrs_0_sepc),
    .csrs_0_mtval(csr_csrs_0_mtval),
    .csrs_0_stval(csr_csrs_0_stval),
    .csrs_0_mtvec(csr_csrs_0_mtvec),
    .csrs_0_stvec(csr_csrs_0_stvec),
    .csrs_0_mcause(csr_csrs_0_mcause),
    .csrs_0_scause(csr_csrs_0_scause),
    .csrs_0_satp(csr_csrs_0_satp),
    .csrs_0_mip(csr_csrs_0_mip),
    .csrs_0_mie(csr_csrs_0_mie),
    .csrs_0_mscratch(csr_csrs_0_mscratch),
    .csrs_0_sscratch(csr_csrs_0_sscratch),
    .csrs_0_mideleg(csr_csrs_0_mideleg),
    .csrs_0_medeleg(csr_csrs_0_medeleg),
    .current_mode_0(csr_current_mode_0),
    .REG_0(csr_REG_0)
  );
  assign io_fb_bmfs_redirect_kill = wbReBranch | csr_io_event_io_except_kill; // @[Backend.scala 488:42]
  assign io_fb_bmfs_redirect_pc = _io_fb_bmfs_redirect_pc_T[31:0]; // @[Backend.scala 489:28]
  assign io_fb_bmfs_bpu_v = wbBpuV; // @[Backend.scala 490:30]
  assign io_fb_bmfs_bpu_errpr = wbBpuErrpr; // @[Backend.scala 491:30]
  assign io_fb_bmfs_bpu_pc_br = {{32'd0}, wbBpuPCBr}; // @[Backend.scala 492:30]
  assign io_fb_bmfs_bpu_target = wbBpuTarget; // @[Backend.scala 493:30]
  assign io_fb_bmfs_bpu_taken = wbBpuTaken; // @[Backend.scala 494:30]
  assign io_fb_fmbs_please_wait = ~issueQueue_io_sufficient; // @[Backend.scala 153:29]
  assign io_dcache_req_valid = exMemRealValid | dcacheStall; // @[Backend.scala 312:41]
  assign io_dcache_req_bits_addr = ldstAddr[31:0]; // @[Backend.scala 339:22 Backend.scala 344:18]
  assign io_dcache_req_bits_wdata = exFwdRtData_2; // @[Backend.scala 339:22 Backend.scala 343:18]
  assign io_dcache_req_bits_wen = ~exInsts_2_write_dest; // @[Backend.scala 345:43]
  assign io_dcache_req_bits_mtype = {{1'd0}, _exMemReq_memReq_mtype_T_13}; // @[Backend.scala 339:22 Backend.scala 342:18]
  assign csrs_mstatus = csr_csrs_0_mstatus;
  assign csrs_sstatus = csr_csrs_0_sstatus;
  assign csrs_mepc = csr_csrs_0_mepc;
  assign csrs_sepc = csr_csrs_0_sepc;
  assign csrs_mtval = csr_csrs_0_mtval;
  assign csrs_stval = csr_csrs_0_stval;
  assign csrs_mtvec = csr_csrs_0_mtvec;
  assign csrs_stvec = csr_csrs_0_stvec;
  assign csrs_mcause = csr_csrs_0_mcause;
  assign csrs_scause = csr_csrs_0_scause;
  assign csrs_satp = csr_csrs_0_satp;
  assign csrs_mip = csr_csrs_0_mip;
  assign csrs_mie = csr_csrs_0_mie;
  assign csrs_mscratch = csr_csrs_0_mscratch;
  assign csrs_sscratch = csr_csrs_0_sscratch;
  assign csrs_mideleg = csr_csrs_0_mideleg;
  assign csrs_medeleg = csr_csrs_0_medeleg;
  assign istall_0 = istall;
  assign _WIRE_4_0_0 = nop_ysyx_print;
  assign _WIRE_4_0_1 = nop_ysyx_print;
  assign _WIRE_4_0_2 = _WIRE_4_2;
  assign _WIRE_1_0_0 = _WIRE_1_0;
  assign _WIRE_1_0_1 = _WIRE_1_1;
  assign _WIRE_1_0_2 = _WIRE_1_2;
  assign current_mode = csr_current_mode_0;
  assign _WIRE_0_0 = regFile__WIRE_0_0;
  assign _WIRE_0_1 = regFile__WIRE_0_1;
  assign _WIRE_0_2 = regFile__WIRE_0_2;
  assign _WIRE_0_3 = regFile__WIRE_0_3;
  assign _WIRE_0_4 = regFile__WIRE_0_4;
  assign _WIRE_0_5 = regFile__WIRE_0_5;
  assign _WIRE_0_6 = regFile__WIRE_0_6;
  assign _WIRE_0_7 = regFile__WIRE_0_7;
  assign _WIRE_0_8 = regFile__WIRE_0_8;
  assign _WIRE_0_9 = regFile__WIRE_0_9;
  assign _WIRE_0_10 = regFile__WIRE_0_10;
  assign _WIRE_0_11 = regFile__WIRE_0_11;
  assign _WIRE_0_12 = regFile__WIRE_0_12;
  assign _WIRE_0_13 = regFile__WIRE_0_13;
  assign _WIRE_0_14 = regFile__WIRE_0_14;
  assign _WIRE_0_15 = regFile__WIRE_0_15;
  assign _WIRE_0_16 = regFile__WIRE_0_16;
  assign _WIRE_0_17 = regFile__WIRE_0_17;
  assign _WIRE_0_18 = regFile__WIRE_0_18;
  assign _WIRE_0_19 = regFile__WIRE_0_19;
  assign _WIRE_0_20 = regFile__WIRE_0_20;
  assign _WIRE_0_21 = regFile__WIRE_0_21;
  assign _WIRE_0_22 = regFile__WIRE_0_22;
  assign _WIRE_0_23 = regFile__WIRE_0_23;
  assign _WIRE_0_24 = regFile__WIRE_0_24;
  assign _WIRE_0_25 = regFile__WIRE_0_25;
  assign _WIRE_0_26 = regFile__WIRE_0_26;
  assign _WIRE_0_27 = regFile__WIRE_0_27;
  assign _WIRE_0_28 = regFile__WIRE_0_28;
  assign _WIRE_0_29 = regFile__WIRE_0_29;
  assign _WIRE_0_30 = regFile__WIRE_0_30;
  assign _WIRE_0_31 = regFile__WIRE_0_31;
  assign dstall_0 = dstall;
  assign _WIRE_6_0 = _WIRE__0;
  assign _WIRE_6_1 = _WIRE__1;
  assign _WIRE_6_2 = _WIRE__2;
  assign counter_0 = counter;
  assign mduStall_0 = mduStall;
  assign _WIRE_3_0_0 = _WIRE_3_0;
  assign _WIRE_3_0_1 = _WIRE_3_1;
  assign _WIRE_3_0_2 = _WIRE_3_2;
  assign common_0 = common;
  assign _WIRE_5_0_0 = _WIRE_5_0;
  assign _WIRE_5_0_1 = _WIRE_5_1;
  assign _WIRE_5_0_2 = _WIRE_5_2;
  assign instret_0 = instret;
  assign _WIRE_2_0_0 = _WIRE_2_0;
  assign _WIRE_2_0_1 = _WIRE_2_1;
  assign _WIRE_2_0_2 = _WIRE_2_2;
  assign REG_0 = csr_REG_0;
  assign wbInsts_0_ysyx_debug = wbInsts__0_ysyx_debug;
  assign alu_io_a = 2'h1 == exInsts_0_src_a ? _alu_io_a_T : _alu_io_a_T_2; // @[Mux.scala 80:57]
  assign alu_io_b = exInsts_0_src_b == 2'h0 ? exFwdRtData_0 : genImm_0; // @[Backend.scala 289:18]
  assign alu_io_aluOp = exInsts_0_alu_op; // @[Backend.scala 290:16]
  assign alu_io_aluExpand = exInsts_0_alu_expand; // @[Backend.scala 291:20]
  assign alu_io_aluCsr = exInsts_0_src_b == 2'h2; // @[Backend.scala 292:37]
  assign alu_io_csr = csr_io_common_io_out; // @[Backend.scala 293:14]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_kill = io_fb_bmfs_redirect_kill; // @[Backend.scala 303:15]
  assign mdu_io_req_valid = exInstsValid_1 & _aluValid_T; // @[Backend.scala 280:33]
  assign mdu_io_req_op = exInsts_1_alu_op; // @[Backend.scala 301:17]
  assign mdu_io_req_expand = exInsts_1_alu_expand; // @[Backend.scala 302:21]
  assign mdu_io_req_in1 = exInsts_1_src_a == 2'h0 ? exFwdRsData_1 : {{32'd0}, exInsts_1_pc}; // @[Backend.scala 299:24]
  assign mdu_io_req_in2 = exInsts_1_src_b == 2'h0 ? exFwdRtData_1 : genImm_1; // @[Backend.scala 300:24]
  assign issueQueue_clock = clock;
  assign issueQueue_reset = reset;
  assign issueQueue_io_enqStep = {{2'd0}, io_fb_fmbs_instn}; // @[Backend.scala 158:25]
  assign issueQueue_io_enqReq = io_fb_fmbs_instn != 2'h0; // @[Backend.scala 157:45]
  assign issueQueue_io_deqStep = {{2'd0}, issueArbiter_io_issue_num}; // @[Backend.scala 64:26 Backend.scala 171:31]
  assign issueQueue_io_deqReq = ~bubble_w & ~(|issueQueue_io_items & issueNum == 2'h0); // @[Backend.scala 156:37]
  assign issueQueue_io_din_0_illegal = io_fb_fmbs_inst_ops_0[160]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_next_pc = io_fb_fmbs_inst_ops_0[159:156]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_alu_mdu_lsu = io_fb_fmbs_inst_ops_0[155:154]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_branch_type = io_fb_fmbs_inst_ops_0[153:150]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_src_a = io_fb_fmbs_inst_ops_0[149:148]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_src_b = io_fb_fmbs_inst_ops_0[147:146]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_write_dest = io_fb_fmbs_inst_ops_0[145]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_alu_op = io_fb_fmbs_inst_ops_0[144:140]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_alu_expand = io_fb_fmbs_inst_ops_0[139]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_mem_width = io_fb_fmbs_inst_ops_0[138:136]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_write_src = io_fb_fmbs_inst_ops_0[135:134]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_rs1 = io_fb_fmbs_inst_ops_0[133:129]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_rs2 = io_fb_fmbs_inst_ops_0[128:124]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_rd = io_fb_fmbs_inst_ops_0[123:119]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_imm = io_fb_fmbs_inst_ops_0[118:99]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_pc = io_fb_fmbs_inst_ops_0[98:67]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_predict_taken = io_fb_fmbs_inst_ops_0[66]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_target_pc = io_fb_fmbs_inst_ops_0[65:34]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_ysyx_debug = io_fb_fmbs_inst_ops_0[33]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_ysyx_print = io_fb_fmbs_inst_ops_0[32]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_0_inst = io_fb_fmbs_inst_ops_0[31:0]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_illegal = io_fb_fmbs_inst_ops_1[160]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_next_pc = io_fb_fmbs_inst_ops_1[159:156]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_alu_mdu_lsu = io_fb_fmbs_inst_ops_1[155:154]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_branch_type = io_fb_fmbs_inst_ops_1[153:150]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_src_a = io_fb_fmbs_inst_ops_1[149:148]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_src_b = io_fb_fmbs_inst_ops_1[147:146]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_write_dest = io_fb_fmbs_inst_ops_1[145]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_alu_op = io_fb_fmbs_inst_ops_1[144:140]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_alu_expand = io_fb_fmbs_inst_ops_1[139]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_mem_width = io_fb_fmbs_inst_ops_1[138:136]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_write_src = io_fb_fmbs_inst_ops_1[135:134]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_rs1 = io_fb_fmbs_inst_ops_1[133:129]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_rs2 = io_fb_fmbs_inst_ops_1[128:124]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_rd = io_fb_fmbs_inst_ops_1[123:119]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_imm = io_fb_fmbs_inst_ops_1[118:99]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_pc = io_fb_fmbs_inst_ops_1[98:67]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_predict_taken = io_fb_fmbs_inst_ops_1[66]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_target_pc = io_fb_fmbs_inst_ops_1[65:34]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_ysyx_debug = io_fb_fmbs_inst_ops_1[33]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_ysyx_print = io_fb_fmbs_inst_ops_1[32]; // @[Backend.scala 163:60]
  assign issueQueue_io_din_1_inst = io_fb_fmbs_inst_ops_1[31:0]; // @[Backend.scala 163:60]
  assign issueQueue_io_flush = io_fb_bmfs_redirect_kill; // @[Backend.scala 154:25]
  assign issueArbiter_io_insts_in_0_illegal = issueQueue_io_dout_0_illegal; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_next_pc = issueQueue_io_dout_0_next_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_alu_mdu_lsu = issueQueue_io_dout_0_alu_mdu_lsu; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_branch_type = issueQueue_io_dout_0_branch_type; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_src_a = issueQueue_io_dout_0_src_a; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_src_b = issueQueue_io_dout_0_src_b; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_write_dest = issueQueue_io_dout_0_write_dest; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_alu_op = issueQueue_io_dout_0_alu_op; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_alu_expand = issueQueue_io_dout_0_alu_expand; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_mem_width = issueQueue_io_dout_0_mem_width; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_write_src = issueQueue_io_dout_0_write_src; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_rs1 = issueQueue_io_dout_0_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_rs2 = issueQueue_io_dout_0_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_rd = issueQueue_io_dout_0_rd; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_imm = issueQueue_io_dout_0_imm; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_pc = issueQueue_io_dout_0_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_predict_taken = issueQueue_io_dout_0_predict_taken; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_target_pc = issueQueue_io_dout_0_target_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_ysyx_debug = issueQueue_io_dout_0_ysyx_debug; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_ysyx_print = issueQueue_io_dout_0_ysyx_print; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_0_inst = issueQueue_io_dout_0_inst; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_illegal = issueQueue_io_dout_1_illegal; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_next_pc = issueQueue_io_dout_1_next_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_alu_mdu_lsu = issueQueue_io_dout_1_alu_mdu_lsu; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_branch_type = issueQueue_io_dout_1_branch_type; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_src_a = issueQueue_io_dout_1_src_a; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_src_b = issueQueue_io_dout_1_src_b; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_write_dest = issueQueue_io_dout_1_write_dest; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_alu_op = issueQueue_io_dout_1_alu_op; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_alu_expand = issueQueue_io_dout_1_alu_expand; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_mem_width = issueQueue_io_dout_1_mem_width; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_write_src = issueQueue_io_dout_1_write_src; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_rs1 = issueQueue_io_dout_1_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_rs2 = issueQueue_io_dout_1_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_rd = issueQueue_io_dout_1_rd; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_imm = issueQueue_io_dout_1_imm; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_pc = issueQueue_io_dout_1_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_predict_taken = issueQueue_io_dout_1_predict_taken; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_target_pc = issueQueue_io_dout_1_target_pc; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_ysyx_debug = issueQueue_io_dout_1_ysyx_debug; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_ysyx_print = issueQueue_io_dout_1_ysyx_print; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_insts_in_1_inst = issueQueue_io_dout_1_inst; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign issueArbiter_io_queue_items = issueQueue_io_items; // @[Backend.scala 166:31]
  assign issueArbiter_io_ld_dest_ex = _issueArbiter_io_ld_dest_ex_T_1 & exInsts_2_rd; // @[Backend.scala 167:73]
  assign issueArbiter_io_rss_in_0 = exInstsValid_1 & exInsts_1_write_dest & exInsts_1_rd != 5'h0 ? _GEN_32 : _GEN_28; // @[Backend.scala 205:96]
  assign issueArbiter_io_rss_in_1 = exInstsValid_1 & exInsts_1_write_dest & exInsts_1_rd != 5'h0 ? _GEN_34 : _GEN_30; // @[Backend.scala 205:96]
  assign issueArbiter_io_rts_in_0 = exInstsValid_1 & exInsts_1_write_dest & exInsts_1_rd != 5'h0 ? _GEN_33 : _GEN_29; // @[Backend.scala 205:96]
  assign issueArbiter_io_rts_in_1 = exInstsValid_1 & exInsts_1_write_dest & exInsts_1_rd != 5'h0 ? _GEN_35 : _GEN_31; // @[Backend.scala 205:96]
  assign regFile_clock = clock;
  assign regFile_reset = reset;
  assign regFile_io_rs_addr_vec_0 = issueQueue_io_dout_0_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign regFile_io_rs_addr_vec_1 = issueQueue_io_dout_0_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign regFile_io_rs_addr_vec_2 = issueQueue_io_dout_1_rs1; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign regFile_io_rs_addr_vec_3 = issueQueue_io_dout_1_rs2; // @[Backend.scala 65:26 Backend.scala 160:19]
  assign regFile_io_wen_vec_0 = wbInstsValid_0 ? _regFile_io_wen_vec_0_T_2 : _regFile_io_wen_vec_0_T_6; // @[Backend.scala 497:31]
  assign regFile_io_wen_vec_1 = wbInstsValid_2 ? _regFile_io_wen_vec_1_T_2 : _regFile_io_wen_vec_0_T_6; // @[Backend.scala 504:31]
  assign regFile_io_rd_addr_vec_0 = wbInstsValid_0 ? wbInsts__0_rd : wbInsts__1_rd; // @[Backend.scala 501:35]
  assign regFile_io_rd_addr_vec_1 = wbInstsValid_2 ? wbInsts__2_rd : wbInsts__1_rd; // @[Backend.scala 509:35]
  assign regFile_io_rd_data_vec_0 = wbInstsValid_0 ? wbResult_0 : wbResult_1; // @[Backend.scala 502:35]
  assign regFile_io_rd_data_vec_1 = wbInstsValid_2 ? wbLdData : wbResult_1; // @[Backend.scala 508:35]
  assign regFile_difftestSaddr = difftest_saddr;
  assign regFile_difftestSval = difftest_sval;
  assign regFile_difftestSync = difftest_sync;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_common_io_in = wbCsrData; // @[Backend.scala 572:31]
  assign csr_io_common_io_wen = csrWbValid & wbInstsValid_0; // @[Backend.scala 570:45]
  assign csr_io_common_io_num = csr_io_common_io_wen ? wbInsts__0_imm[11:0] : exInsts_0_imm[11:0]; // @[Backend.scala 571:37]
  assign csr_io_event_io_exception_vec_2 = wbInsts__0_illegal & wbInstsValid_0; // @[Backend.scala 519:42]
  assign csr_io_event_io_exception_vec_3 = wbInsts__0_next_pc == 4'h8 & wbInstsValid_0; // @[Backend.scala 518:64]
  assign csr_io_event_io_exception_vec_4 = wbLdMaReal | wbFetchMaReal; // @[Backend.scala 535:59]
  assign csr_io_event_io_exception_vec_6 = wbInstsValid_2 & wbStMa; // @[Backend.scala 516:39]
  assign csr_io_event_io_deal_with_int = wbInterruptd & |_wb_deal_with_int_T & exInterruptd; // @[Backend.scala 542:91]
  assign csr_io_event_io_is_mret = wbInsts__0_next_pc == 4'h6 & wbInstsValid_0; // @[Backend.scala 557:74]
  assign csr_io_event_io_is_sret = wbInsts__0_next_pc == 4'h7 & wbInstsValid_0; // @[Backend.scala 558:74]
  assign csr_io_event_io_is_ecall = wbInsts__0_next_pc == 4'h5 & wbInstsValid_0; // @[Backend.scala 517:63]
  assign csr_io_event_io_bad_address = {{32'd0}, _csr_io_event_io_bad_address_T}; // @[Backend.scala 567:37]
  assign csr_io_event_io_epc = wb_deal_with_int ? wb_pc_min : {{32'd0}, _csr_io_event_io_epc_T_2}; // @[Backend.scala 565:37]
  always @(posedge clock) begin
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_illegal <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_illegal <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_illegal <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_illegal <= issueArbiter_io_insts_out_0_illegal; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_next_pc <= 4'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_next_pc <= 4'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_next_pc <= 4'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_next_pc <= issueArbiter_io_insts_out_0_next_pc; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_alu_mdu_lsu <= 2'h3; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_alu_mdu_lsu <= 2'h3; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_alu_mdu_lsu <= 2'h3; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_alu_mdu_lsu <= issueArbiter_io_insts_out_0_alu_mdu_lsu; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_branch_type <= 4'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_branch_type <= 4'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_branch_type <= 4'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_branch_type <= issueArbiter_io_insts_out_0_branch_type; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_src_a <= 2'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_src_a <= 2'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_src_a <= 2'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_src_a <= issueArbiter_io_insts_out_0_src_a; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_src_b <= 2'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_src_b <= 2'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_src_b <= 2'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_src_b <= issueArbiter_io_insts_out_0_src_b; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_write_dest <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_write_dest <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_write_dest <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_write_dest <= issueArbiter_io_insts_out_0_write_dest; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_alu_op <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_alu_op <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_alu_op <= 5'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_alu_op <= issueArbiter_io_insts_out_0_alu_op; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_alu_expand <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_alu_expand <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_alu_expand <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_alu_expand <= issueArbiter_io_insts_out_0_alu_expand; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_write_src <= 2'h1; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_write_src <= 2'h1; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_write_src <= 2'h1; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_write_src <= issueArbiter_io_insts_out_0_write_src; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_rs1 <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_rs1 <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_rs1 <= 5'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_rs1 <= issueArbiter_io_insts_out_0_rs1; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_rd <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_rd <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_rd <= 5'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_rd <= issueArbiter_io_insts_out_0_rd; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_imm <= 20'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_imm <= 20'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_imm <= 20'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_imm <= issueArbiter_io_insts_out_0_imm; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_pc <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_pc <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_pc <= issueInsts_0_pc; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_pc <= issueArbiter_io_insts_out_0_pc; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_predict_taken <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_predict_taken <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_predict_taken <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_predict_taken <= issueArbiter_io_insts_out_0_predict_taken; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_target_pc <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_target_pc <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_target_pc <= 32'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_target_pc <= issueArbiter_io_insts_out_0_target_pc; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_ysyx_debug <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_ysyx_debug <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_ysyx_debug <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_ysyx_debug <= issueArbiter_io_insts_out_0_ysyx_debug; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_ysyx_print <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_ysyx_print <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_ysyx_print <= 1'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_ysyx_print <= issueArbiter_io_insts_out_0_ysyx_print; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_0_inst <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_0_inst <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInsts_0_inst <= 32'h0; // @[Backend.scala 257:18]
      end else begin
        exInsts_0_inst <= issueArbiter_io_insts_out_0_inst; // @[Backend.scala 263:20]
      end
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_src_a <= 2'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_src_a <= 2'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_src_a <= issueArbiter_io_insts_out_1_src_a; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_src_b <= 2'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_src_b <= 2'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_src_b <= issueArbiter_io_insts_out_1_src_b; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_write_dest <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_write_dest <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_write_dest <= issueArbiter_io_insts_out_1_write_dest; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_alu_op <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_alu_op <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_alu_op <= issueArbiter_io_insts_out_1_alu_op; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_alu_expand <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_alu_expand <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_alu_expand <= issueArbiter_io_insts_out_1_alu_expand; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_rd <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_rd <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_rd <= issueArbiter_io_insts_out_1_rd; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_imm <= 20'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_imm <= 20'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_imm <= issueArbiter_io_insts_out_1_imm; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_pc <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_pc <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_pc <= issueArbiter_io_insts_out_1_pc; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_ysyx_print <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_ysyx_print <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_ysyx_print <= issueArbiter_io_insts_out_1_ysyx_print; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_1_inst <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_1_inst <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_1_inst <= issueArbiter_io_insts_out_1_inst; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_src_a <= 2'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_src_a <= 2'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_src_a <= issueArbiter_io_insts_out_2_src_a; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_write_dest <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_write_dest <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_write_dest <= issueArbiter_io_insts_out_2_write_dest; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_alu_op <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_alu_op <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_alu_op <= issueArbiter_io_insts_out_2_alu_op; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_mem_width <= 3'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_mem_width <= 3'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_mem_width <= issueArbiter_io_insts_out_2_mem_width; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_rd <= 5'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_rd <= 5'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_rd <= issueArbiter_io_insts_out_2_rd; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_imm <= 20'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_imm <= 20'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_imm <= issueArbiter_io_insts_out_2_imm; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_pc <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_pc <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_pc <= issueArbiter_io_insts_out_2_pc; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_ysyx_print <= 1'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_ysyx_print <= 1'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_ysyx_print <= issueArbiter_io_insts_out_2_ysyx_print; // @[Backend.scala 266:18]
    end
    if (reset) begin // @[Backend.scala 81:29]
      exInsts_2_inst <= 32'h0; // @[Backend.scala 81:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInsts_2_inst <= 32'h0; // @[Backend.scala 248:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInsts_2_inst <= issueArbiter_io_insts_out_2_inst; // @[Backend.scala 266:18]
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 245:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
        exInstsOrder_0 <= issueArbiter_io_insts_order_0; // @[Backend.scala 252:18]
      end
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 245:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
        exInstsOrder_1 <= issueArbiter_io_insts_order_1; // @[Backend.scala 252:18]
      end
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 245:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
        exInstsOrder_2 <= issueArbiter_io_insts_order_2; // @[Backend.scala 252:18]
      end
    end
    if (reset) begin // @[Backend.scala 83:29]
      exInstsValid_0 <= 1'h0; // @[Backend.scala 83:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInstsValid_0 <= 1'h0; // @[Backend.scala 249:23]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInstsValid_0 <= |_exInstsValid_0_T; // @[Backend.scala 254:23]
      end else begin
        exInstsValid_0 <= issueArbiter_io_issue_fu_valid_0; // @[Backend.scala 262:20]
      end
    end
    if (reset) begin // @[Backend.scala 83:29]
      exInstsValid_1 <= 1'h0; // @[Backend.scala 83:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInstsValid_1 <= 1'h0; // @[Backend.scala 249:23]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInstsValid_1 <= 1'h0; // @[Backend.scala 259:25]
      end else begin
        exInstsValid_1 <= issueArbiter_io_issue_fu_valid_1; // @[Backend.scala 262:20]
      end
    end
    if (reset) begin // @[Backend.scala 83:29]
      exInstsValid_2 <= 1'h0; // @[Backend.scala 83:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInstsValid_2 <= 1'h0; // @[Backend.scala 249:23]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      if (csr_io_event_io_call_for_int) begin // @[Backend.scala 253:41]
        exInstsValid_2 <= 1'h0; // @[Backend.scala 259:25]
      end else begin
        exInstsValid_2 <= issueArbiter_io_issue_fu_valid_2; // @[Backend.scala 262:20]
      end
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRsData_0 <= issueRss_0; // @[Backend.scala 273:22]
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRsData_1 <= issueRss_1; // @[Backend.scala 273:22]
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRsData_2 <= issueRss_2; // @[Backend.scala 273:22]
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRtData_0 <= issueRts_0; // @[Backend.scala 274:22]
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRtData_1 <= issueRts_1; // @[Backend.scala 274:22]
    end
    if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 271:19]
      exFwdRtData_2 <= issueRts_2; // @[Backend.scala 274:22]
    end
    if (reset) begin // @[Backend.scala 99:29]
      exInterruptd <= 1'h0; // @[Backend.scala 99:29]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 245:17]
      exInterruptd <= 1'h0; // @[Backend.scala 246:18]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 251:24]
      exInterruptd <= csr_io_event_io_call_for_int; // @[Backend.scala 268:18]
    end
    reBranchPC <= _GEN_386[31:0];
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        if (exInsts_0_write_src == 2'h3 | exInsts_0_next_pc != 4'h0) begin // @[Backend.scala 423:19]
          wbResult_0 <= {{32'd0}, _exReBranchPC_T_3};
        end else if (2'h2 == exInsts_0_src_b) begin // @[Mux.scala 80:57]
          wbResult_0 <= csr_io_common_io_out;
        end else begin
          wbResult_0 <= alu_io_r;
        end
      end
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbResult_1 <= mdu_io_resp_r; // @[Backend.scala 474:17]
      end
    end
    if (reset) begin // @[Backend.scala 126:33]
      wbInstsValid_0 <= 1'h0; // @[Backend.scala 126:33]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 455:17]
      wbInstsValid_0 <= 1'h0; // @[Backend.scala 457:23]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
      wbInstsValid_0 <= exInstsTrueValid_0; // @[Backend.scala 469:23]
    end
    if (reset) begin // @[Backend.scala 126:33]
      wbInstsValid_1 <= 1'h0; // @[Backend.scala 126:33]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 455:17]
      wbInstsValid_1 <= 1'h0; // @[Backend.scala 457:23]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
      wbInstsValid_1 <= exInstsTrueValid_1; // @[Backend.scala 469:23]
    end
    if (reset) begin // @[Backend.scala 126:33]
      wbInstsValid_2 <= 1'h0; // @[Backend.scala 126:33]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 455:17]
      wbInstsValid_2 <= dcacheStall; // @[Backend.scala 459:21]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
      wbInstsValid_2 <= ldstValid; // @[Backend.scala 469:23]
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInstsOrder_0 <= exInstsOrder_0; // @[Backend.scala 472:18]
      end
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInstsOrder_1 <= exInstsOrder_1; // @[Backend.scala 472:18]
      end
    end
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInstsOrder_2 <= exInstsOrder_2; // @[Backend.scala 472:18]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_illegal <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_illegal <= exInsts_0_illegal; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_next_pc <= 4'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_next_pc <= exInsts_0_next_pc; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_alu_mdu_lsu <= 2'h3; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_alu_mdu_lsu <= exInsts_0_alu_mdu_lsu; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_write_dest <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_write_dest <= exInsts_0_write_dest; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_rd <= 5'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_rd <= exInsts_0_rd; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_imm <= 20'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_imm <= exInsts_0_imm; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_pc <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_pc <= exInsts_0_pc; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_ysyx_debug <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_ysyx_debug <= exInsts_0_ysyx_debug; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_ysyx_print <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_ysyx_print <= exInsts_0_ysyx_print; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__0_inst <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__0_inst <= exInsts_0_inst; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__1_write_dest <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__1_write_dest <= exInsts_1_write_dest; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__1_rd <= 5'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__1_rd <= exInsts_1_rd; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__1_pc <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__1_pc <= exInsts_1_pc; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__1_ysyx_print <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__1_ysyx_print <= exInsts_1_ysyx_print; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__1_inst <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__1_inst <= exInsts_1_inst; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_write_dest <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_write_dest <= exInsts_2_write_dest; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_mem_width <= 3'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_mem_width <= exInsts_2_mem_width; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_rd <= 5'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_rd <= exInsts_2_rd; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_pc <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_pc <= exInsts_2_pc; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_ysyx_print <= 1'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_ysyx_print <= exInsts_2_ysyx_print; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 128:33]
      wbInsts__2_inst <= 32'h0; // @[Backend.scala 128:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInsts__2_inst <= exInsts_2_inst; // @[Backend.scala 471:13]
      end
    end
    if (reset) begin // @[Backend.scala 134:33]
      wbReBranch <= 1'h0; // @[Backend.scala 134:33]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 455:17]
      wbReBranch <= 1'h0; // @[Backend.scala 460:16]
    end else if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
      wbReBranch <= reBranch; // @[Backend.scala 481:16]
    end
    wbMisalignedAddr <= io_dcache_req_bits_addr; // @[Backend.scala 137:33]
    if (reset) begin // @[Backend.scala 138:33]
      wbInterruptd <= 1'h0; // @[Backend.scala 138:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbInterruptd <= exInterruptd & _aluValid_T; // @[Backend.scala 463:18]
      end
    end
    if (reset) begin // @[Backend.scala 139:33]
      wbLdMa <= 1'h0; // @[Backend.scala 139:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbLdMa <= ldMisaligned; // @[Backend.scala 475:12]
      end
    end
    if (reset) begin // @[Backend.scala 140:33]
      wbStMa <= 1'h0; // @[Backend.scala 140:33]
    end else if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbStMa <= stMisaligned; // @[Backend.scala 476:12]
      end
    end
    if (reset) begin // @[Backend.scala 141:33]
      wbBpuV <= 1'h0; // @[Backend.scala 141:33]
    end else if (io_fb_bmfs_redirect_kill) begin // @[Backend.scala 455:17]
      wbBpuV <= 1'h0; // @[Backend.scala 461:12]
    end else begin
      wbBpuV <= _GEN_230;
    end
    wbBpuErrpr <= isExPCBr & exInsts_0_target_pc[31:2] != brPC[31:2] & reBranchBrTaken | _bpuErrpr_T_8; // @[Backend.scala 117:114]
    wbBpuPCBr <= {wbBpuPCBr_hi,wbBpuPCBr_lo}; // @[Cat.scala 30:58]
    if (isExPCBr) begin // @[Backend.scala 120:22]
      wbBpuTarget <= brPC;
    end else begin
      wbBpuTarget <= {{32'd0}, jumpPc};
    end
    wbBpuTaken <= reBranchBrTaken | isExPCJump; // @[Backend.scala 121:35]
    if (!(io_fb_bmfs_redirect_kill)) begin // @[Backend.scala 455:17]
      if (_issueQueue_io_deqReq_T) begin // @[Backend.scala 462:26]
        wbCsrData <= alu_io_r; // @[Backend.scala 478:15]
      end
    end
    if (reset) begin // @[Backend.scala 306:30]
      wbMemReqValid <= 1'h0; // @[Backend.scala 306:30]
    end else if (~dcacheStall) begin // @[Backend.scala 349:23]
      wbMemReqValid <= exMemRealValid; // @[Backend.scala 350:19]
    end
    if (reset) begin // @[Backend.scala 315:25]
      wbMemReq_addr <= 32'h0; // @[Backend.scala 315:25]
    end else if (~dcacheStall) begin // @[Backend.scala 349:23]
      wbMemReq_addr <= exMemReq_addr; // @[Backend.scala 351:14]
    end
    if (dcacheStall & ~REG) begin // @[Backend.scala 591:48]
      bufInsts0_pc <= wbInsts__0_pc; // @[Backend.scala 592:17]
    end
    if (dcacheStall & ~REG) begin // @[Backend.scala 591:48]
      bufInsts0_inst <= wbInsts__0_inst; // @[Backend.scala 592:17]
    end
    if (dcacheStall & ~REG) begin // @[Backend.scala 591:48]
      bufInstsValid0 <= wbInstsValid_0; // @[Backend.scala 593:22]
    end
    if (dcacheStall & ~REG) begin // @[Backend.scala 591:48]
      bufInstsOrder0 <= wbInstsOrder_0; // @[Backend.scala 594:22]
    end
    REG <= wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
    tmp_REG <= wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
    if (tmp_REG) begin // @[Backend.scala 598:20]
      REG_1 <= bufInstsValid0 & _issueQueue_io_deqReq_T & |bufInsts0_inst;
    end else begin
      REG_1 <= wbInstsValid_0 & _issueQueue_io_deqReq_T & |wbInsts__0_inst;
    end
    REG_2 <= _tmp_T_13 & _tmp_T_14; // @[Backend.scala 600:49]
    REG_3 <= _tmp_T_21 & _tmp_T_22; // @[Backend.scala 600:49]
    tmp_REG_3 <= wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
    if (tmp_REG_3) begin // @[Backend.scala 603:20]
      if (bufInstsValid0) begin // @[Backend.scala 603:46]
        REG_4 <= bufInsts0_pc;
      end else begin
        REG_4 <= 32'h0;
      end
    end else if (wbInstsValid_0) begin // @[Backend.scala 603:86]
      REG_4 <= wbInsts__0_pc;
    end else begin
      REG_4 <= 32'h0;
    end
    if (wbInstsValid_1) begin // @[Backend.scala 605:23]
      REG_5 <= wbInsts__1_pc;
    end else begin
      REG_5 <= 32'h0;
    end
    if (wbInstsValid_2) begin // @[Backend.scala 605:23]
      REG_6 <= wbInsts__2_pc;
    end else begin
      REG_6 <= 32'h0;
    end
    tmp_REG_6 <= wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
    if (tmp_REG_6) begin // @[Backend.scala 608:20]
      REG_7 <= bufInstsOrder0;
    end else begin
      REG_7 <= wbInstsOrder_0;
    end
    REG_8 <= wbInstsOrder_1; // @[Backend.scala 610:19]
    REG_9 <= wbInstsOrder_2; // @[Backend.scala 610:19]
    tmp_REG_9 <= wbMemReqValid & ~io_dcache_resp_valid; // @[Backend.scala 307:32]
    if (tmp_REG_9) begin // @[Backend.scala 613:20]
      REG_10 <= bufInsts0_inst;
    end else begin
      REG_10 <= wbInsts__0_inst;
    end
    REG_11 <= wbInsts__1_inst; // @[Backend.scala 615:19]
    REG_12 <= wbInsts__2_inst; // @[Backend.scala 615:19]
    REG_13 <= io_dcache_resp_valid & ~wbMemReq_addr[31]; // @[Backend.scala 617:94]
    REG_14 <= wbInsts__0_ysyx_print; // @[Backend.scala 623:60]
    REG_15 <= wbInsts__1_ysyx_print; // @[Backend.scala 623:60]
    REG_16 <= wbInsts__2_ysyx_print; // @[Backend.scala 623:60]
    if (reset) begin // @[Backend.scala 627:26]
      instret <= 64'h0; // @[Backend.scala 627:26]
    end else if (!(bubble_w)) begin // @[Backend.scala 639:19]
      instret <= _instret_T_11;
    end
    if (reset) begin // @[Backend.scala 628:26]
      counter <= 64'h0; // @[Backend.scala 628:26]
    end else begin
      counter <= _counter_T_1; // @[Backend.scala 638:13]
    end
    if (reset) begin // @[Backend.scala 629:25]
      dstall <= 64'h0; // @[Backend.scala 629:25]
    end else begin
      dstall <= _dstall_T_2; // @[Backend.scala 635:12]
    end
    if (reset) begin // @[Backend.scala 631:25]
      istall <= 64'h0; // @[Backend.scala 631:25]
    end else begin
      istall <= _istall_T_2; // @[Backend.scala 636:12]
    end
    if (reset) begin // @[Backend.scala 632:27]
      mduStall <= 64'h0; // @[Backend.scala 632:27]
    end else begin
      mduStall <= _mduStall_T_2; // @[Backend.scala 640:14]
    end
    if (reset) begin // @[Backend.scala 633:25]
      common <= 64'h0; // @[Backend.scala 633:25]
    end else begin
      common <= _common_T_3; // @[Backend.scala 637:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exInsts_0_illegal = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  exInsts_0_next_pc = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  exInsts_0_alu_mdu_lsu = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  exInsts_0_branch_type = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  exInsts_0_src_a = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  exInsts_0_src_b = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  exInsts_0_write_dest = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exInsts_0_alu_op = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  exInsts_0_alu_expand = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exInsts_0_write_src = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  exInsts_0_rs1 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  exInsts_0_rd = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  exInsts_0_imm = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  exInsts_0_pc = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  exInsts_0_predict_taken = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exInsts_0_target_pc = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  exInsts_0_ysyx_debug = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  exInsts_0_ysyx_print = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exInsts_0_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  exInsts_1_src_a = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  exInsts_1_src_b = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  exInsts_1_write_dest = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exInsts_1_alu_op = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  exInsts_1_alu_expand = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  exInsts_1_rd = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  exInsts_1_imm = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  exInsts_1_pc = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  exInsts_1_ysyx_print = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  exInsts_1_inst = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  exInsts_2_src_a = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  exInsts_2_write_dest = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  exInsts_2_alu_op = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  exInsts_2_mem_width = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  exInsts_2_rd = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  exInsts_2_imm = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  exInsts_2_pc = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  exInsts_2_ysyx_print = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  exInsts_2_inst = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  exInstsOrder_0 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  exInstsOrder_1 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  exInstsOrder_2 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  exInstsValid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  exInstsValid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  exInstsValid_2 = _RAND_43[0:0];
  _RAND_44 = {2{`RANDOM}};
  exFwdRsData_0 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  exFwdRsData_1 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  exFwdRsData_2 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  exFwdRtData_0 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  exFwdRtData_1 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  exFwdRtData_2 = _RAND_49[63:0];
  _RAND_50 = {1{`RANDOM}};
  exInterruptd = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  reBranchPC = _RAND_51[31:0];
  _RAND_52 = {2{`RANDOM}};
  wbResult_0 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  wbResult_1 = _RAND_53[63:0];
  _RAND_54 = {1{`RANDOM}};
  wbInstsValid_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  wbInstsValid_1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  wbInstsValid_2 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  wbInstsOrder_0 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  wbInstsOrder_1 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  wbInstsOrder_2 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  wbInsts__0_illegal = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  wbInsts__0_next_pc = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  wbInsts__0_alu_mdu_lsu = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  wbInsts__0_write_dest = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  wbInsts__0_rd = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  wbInsts__0_imm = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  wbInsts__0_pc = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  wbInsts__0_ysyx_debug = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  wbInsts__0_ysyx_print = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  wbInsts__0_inst = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  wbInsts__1_write_dest = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  wbInsts__1_rd = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  wbInsts__1_pc = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  wbInsts__1_ysyx_print = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  wbInsts__1_inst = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  wbInsts__2_write_dest = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  wbInsts__2_mem_width = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  wbInsts__2_rd = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  wbInsts__2_pc = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  wbInsts__2_ysyx_print = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  wbInsts__2_inst = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  wbReBranch = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  wbMisalignedAddr = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  wbInterruptd = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  wbLdMa = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  wbStMa = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  wbBpuV = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  wbBpuErrpr = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  wbBpuPCBr = _RAND_88[31:0];
  _RAND_89 = {2{`RANDOM}};
  wbBpuTarget = _RAND_89[63:0];
  _RAND_90 = {1{`RANDOM}};
  wbBpuTaken = _RAND_90[0:0];
  _RAND_91 = {2{`RANDOM}};
  wbCsrData = _RAND_91[63:0];
  _RAND_92 = {1{`RANDOM}};
  wbMemReqValid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  wbMemReq_addr = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  bufInsts0_pc = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  bufInsts0_inst = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  bufInstsValid0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  bufInstsOrder0 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  REG = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  tmp_REG = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG_1 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG_2 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG_3 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  tmp_REG_3 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_4 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  REG_5 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  REG_6 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  tmp_REG_6 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_7 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  REG_8 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  REG_9 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  tmp_REG_9 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG_10 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  REG_11 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  REG_12 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  REG_13 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG_14 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_15 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG_16 = _RAND_118[0:0];
  _RAND_119 = {2{`RANDOM}};
  instret = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  counter = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  dstall = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  istall = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  mduStall = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  common = _RAND_124[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  output [31:0] io_icache_req_bits_addr,
  output [2:0]  io_icache_req_bits_mtype,
  input         io_icache_resp_valid,
  input  [31:0] io_icache_resp_bits_rdata_0,
  input  [31:0] io_icache_resp_bits_rdata_1,
  input         io_icache_resp_bits_respn,
  output        io_dcache_req_valid,
  output [31:0] io_dcache_req_bits_addr,
  output [63:0] io_dcache_req_bits_wdata,
  output        io_dcache_req_bits_wen,
  output [2:0]  io_dcache_req_bits_mtype,
  input         io_dcache_resp_valid,
  input  [31:0] io_dcache_resp_bits_rdata_0,
  input  [31:0] io_dcache_resp_bits_rdata_1,
  output [63:0] csrs_mstatus,
  output [63:0] csrs_sstatus,
  output [63:0] csrs_mepc,
  output [63:0] csrs_sepc,
  output [63:0] csrs_mtval,
  output [63:0] csrs_stval,
  output [63:0] csrs_mtvec,
  output [63:0] csrs_stvec,
  output [63:0] csrs_mcause,
  output [63:0] csrs_scause,
  output [63:0] csrs_satp,
  output [63:0] csrs_mip,
  output [63:0] csrs_mie,
  output [63:0] csrs_mscratch,
  output [63:0] csrs_sscratch,
  output [63:0] csrs_mideleg,
  output [63:0] csrs_medeleg,
  output [63:0] istall,
  output        _WIRE_4_0,
  output        _WIRE_4_1,
  output        _WIRE_4_2,
  output [31:0] _WIRE_1_0,
  output [31:0] _WIRE_1_1,
  output [31:0] _WIRE_1_2,
  input  [4:0]  difftest_saddr,
  output [1:0]  current_mode,
  output [63:0] _WIRE__0,
  output [63:0] _WIRE__1,
  output [63:0] _WIRE__2,
  output [63:0] _WIRE__3,
  output [63:0] _WIRE__4,
  output [63:0] _WIRE__5,
  output [63:0] _WIRE__6,
  output [63:0] _WIRE__7,
  output [63:0] _WIRE__8,
  output [63:0] _WIRE__9,
  output [63:0] _WIRE__10,
  output [63:0] _WIRE__11,
  output [63:0] _WIRE__12,
  output [63:0] _WIRE__13,
  output [63:0] _WIRE__14,
  output [63:0] _WIRE__15,
  output [63:0] _WIRE__16,
  output [63:0] _WIRE__17,
  output [63:0] _WIRE__18,
  output [63:0] _WIRE__19,
  output [63:0] _WIRE__20,
  output [63:0] _WIRE__21,
  output [63:0] _WIRE__22,
  output [63:0] _WIRE__23,
  output [63:0] _WIRE__24,
  output [63:0] _WIRE__25,
  output [63:0] _WIRE__26,
  output [63:0] _WIRE__27,
  output [63:0] _WIRE__28,
  output [63:0] _WIRE__29,
  output [63:0] _WIRE__30,
  output [63:0] _WIRE__31,
  output [63:0] dstall,
  output        _WIRE_0_0,
  output        _WIRE_0_1,
  output        _WIRE_0_2,
  output [63:0] counter,
  input  [31:0] difftest_sval,
  output [63:0] mduStall,
  output [31:0] _WIRE_3_0,
  output [31:0] _WIRE_3_1,
  output [31:0] _WIRE_3_2,
  output [63:0] common,
  output        _WIRE_5_0,
  output        _WIRE_5_1,
  output        _WIRE_5_2,
  output [63:0] instret,
  output [1:0]  _WIRE_2_0,
  output [1:0]  _WIRE_2_1,
  output [1:0]  _WIRE_2_2,
  output        REG_0,
  input         difftest_sync,
  output        wbInsts_0_ysyx_debug
);
  wire  fe_clock; // @[Core.scala 97:18]
  wire  fe_reset; // @[Core.scala 97:18]
  wire  fe_io_fb_bmfs_redirect_kill; // @[Core.scala 97:18]
  wire [31:0] fe_io_fb_bmfs_redirect_pc; // @[Core.scala 97:18]
  wire  fe_io_fb_bmfs_bpu_v; // @[Core.scala 97:18]
  wire  fe_io_fb_bmfs_bpu_errpr; // @[Core.scala 97:18]
  wire [63:0] fe_io_fb_bmfs_bpu_pc_br; // @[Core.scala 97:18]
  wire [63:0] fe_io_fb_bmfs_bpu_target; // @[Core.scala 97:18]
  wire  fe_io_fb_bmfs_bpu_taken; // @[Core.scala 97:18]
  wire [1:0] fe_io_fb_fmbs_instn; // @[Core.scala 97:18]
  wire [160:0] fe_io_fb_fmbs_inst_ops_0; // @[Core.scala 97:18]
  wire [160:0] fe_io_fb_fmbs_inst_ops_1; // @[Core.scala 97:18]
  wire  fe_io_fb_fmbs_please_wait; // @[Core.scala 97:18]
  wire  fe_io_icache_req_valid; // @[Core.scala 97:18]
  wire [31:0] fe_io_icache_req_bits_addr; // @[Core.scala 97:18]
  wire [2:0] fe_io_icache_req_bits_mtype; // @[Core.scala 97:18]
  wire  fe_io_icache_resp_valid; // @[Core.scala 97:18]
  wire [31:0] fe_io_icache_resp_bits_rdata_0; // @[Core.scala 97:18]
  wire [31:0] fe_io_icache_resp_bits_rdata_1; // @[Core.scala 97:18]
  wire  fe_io_icache_resp_bits_respn; // @[Core.scala 97:18]
  wire  fe_cache_stall_0; // @[Core.scala 97:18]
  wire  be_clock; // @[Core.scala 98:18]
  wire  be_reset; // @[Core.scala 98:18]
  wire  be_io_fb_bmfs_redirect_kill; // @[Core.scala 98:18]
  wire [31:0] be_io_fb_bmfs_redirect_pc; // @[Core.scala 98:18]
  wire  be_io_fb_bmfs_bpu_v; // @[Core.scala 98:18]
  wire  be_io_fb_bmfs_bpu_errpr; // @[Core.scala 98:18]
  wire [63:0] be_io_fb_bmfs_bpu_pc_br; // @[Core.scala 98:18]
  wire [63:0] be_io_fb_bmfs_bpu_target; // @[Core.scala 98:18]
  wire  be_io_fb_bmfs_bpu_taken; // @[Core.scala 98:18]
  wire [1:0] be_io_fb_fmbs_instn; // @[Core.scala 98:18]
  wire [160:0] be_io_fb_fmbs_inst_ops_0; // @[Core.scala 98:18]
  wire [160:0] be_io_fb_fmbs_inst_ops_1; // @[Core.scala 98:18]
  wire  be_io_fb_fmbs_please_wait; // @[Core.scala 98:18]
  wire  be_io_dcache_req_valid; // @[Core.scala 98:18]
  wire [31:0] be_io_dcache_req_bits_addr; // @[Core.scala 98:18]
  wire [63:0] be_io_dcache_req_bits_wdata; // @[Core.scala 98:18]
  wire  be_io_dcache_req_bits_wen; // @[Core.scala 98:18]
  wire [2:0] be_io_dcache_req_bits_mtype; // @[Core.scala 98:18]
  wire  be_io_dcache_resp_valid; // @[Core.scala 98:18]
  wire [31:0] be_io_dcache_resp_bits_rdata_0; // @[Core.scala 98:18]
  wire [31:0] be_io_dcache_resp_bits_rdata_1; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mstatus; // @[Core.scala 98:18]
  wire [63:0] be_csrs_sstatus; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mepc; // @[Core.scala 98:18]
  wire [63:0] be_csrs_sepc; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mtval; // @[Core.scala 98:18]
  wire [63:0] be_csrs_stval; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mtvec; // @[Core.scala 98:18]
  wire [63:0] be_csrs_stvec; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mcause; // @[Core.scala 98:18]
  wire [63:0] be_csrs_scause; // @[Core.scala 98:18]
  wire [63:0] be_csrs_satp; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mip; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mie; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mscratch; // @[Core.scala 98:18]
  wire [63:0] be_csrs_sscratch; // @[Core.scala 98:18]
  wire [63:0] be_csrs_mideleg; // @[Core.scala 98:18]
  wire [63:0] be_csrs_medeleg; // @[Core.scala 98:18]
  wire [63:0] be_istall_0; // @[Core.scala 98:18]
  wire  be__WIRE_4_0_0; // @[Core.scala 98:18]
  wire  be__WIRE_4_0_1; // @[Core.scala 98:18]
  wire  be__WIRE_4_0_2; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_1_0_0; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_1_0_1; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_1_0_2; // @[Core.scala 98:18]
  wire [4:0] be_difftest_saddr; // @[Core.scala 98:18]
  wire [1:0] be_current_mode; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_0; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_1; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_2; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_3; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_4; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_5; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_6; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_7; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_8; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_9; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_10; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_11; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_12; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_13; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_14; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_15; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_16; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_17; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_18; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_19; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_20; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_21; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_22; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_23; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_24; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_25; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_26; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_27; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_28; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_29; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_30; // @[Core.scala 98:18]
  wire [63:0] be__WIRE_0_31; // @[Core.scala 98:18]
  wire [63:0] be_dstall_0; // @[Core.scala 98:18]
  wire  be__WIRE_6_0; // @[Core.scala 98:18]
  wire  be__WIRE_6_1; // @[Core.scala 98:18]
  wire  be__WIRE_6_2; // @[Core.scala 98:18]
  wire [63:0] be_counter_0; // @[Core.scala 98:18]
  wire  be_icache_stall; // @[Core.scala 98:18]
  wire [31:0] be_difftest_sval; // @[Core.scala 98:18]
  wire [63:0] be_mduStall_0; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_3_0_0; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_3_0_1; // @[Core.scala 98:18]
  wire [31:0] be__WIRE_3_0_2; // @[Core.scala 98:18]
  wire [63:0] be_common_0; // @[Core.scala 98:18]
  wire  be__WIRE_5_0_0; // @[Core.scala 98:18]
  wire  be__WIRE_5_0_1; // @[Core.scala 98:18]
  wire  be__WIRE_5_0_2; // @[Core.scala 98:18]
  wire [63:0] be_instret_0; // @[Core.scala 98:18]
  wire [1:0] be__WIRE_2_0_0; // @[Core.scala 98:18]
  wire [1:0] be__WIRE_2_0_1; // @[Core.scala 98:18]
  wire [1:0] be__WIRE_2_0_2; // @[Core.scala 98:18]
  wire  be_REG_0; // @[Core.scala 98:18]
  wire  be_difftest_sync; // @[Core.scala 98:18]
  wire  be_wbInsts_0_ysyx_debug; // @[Core.scala 98:18]
  Frontend fe ( // @[Core.scala 97:18]
    .clock(fe_clock),
    .reset(fe_reset),
    .io_fb_bmfs_redirect_kill(fe_io_fb_bmfs_redirect_kill),
    .io_fb_bmfs_redirect_pc(fe_io_fb_bmfs_redirect_pc),
    .io_fb_bmfs_bpu_v(fe_io_fb_bmfs_bpu_v),
    .io_fb_bmfs_bpu_errpr(fe_io_fb_bmfs_bpu_errpr),
    .io_fb_bmfs_bpu_pc_br(fe_io_fb_bmfs_bpu_pc_br),
    .io_fb_bmfs_bpu_target(fe_io_fb_bmfs_bpu_target),
    .io_fb_bmfs_bpu_taken(fe_io_fb_bmfs_bpu_taken),
    .io_fb_fmbs_instn(fe_io_fb_fmbs_instn),
    .io_fb_fmbs_inst_ops_0(fe_io_fb_fmbs_inst_ops_0),
    .io_fb_fmbs_inst_ops_1(fe_io_fb_fmbs_inst_ops_1),
    .io_fb_fmbs_please_wait(fe_io_fb_fmbs_please_wait),
    .io_icache_req_valid(fe_io_icache_req_valid),
    .io_icache_req_bits_addr(fe_io_icache_req_bits_addr),
    .io_icache_req_bits_mtype(fe_io_icache_req_bits_mtype),
    .io_icache_resp_valid(fe_io_icache_resp_valid),
    .io_icache_resp_bits_rdata_0(fe_io_icache_resp_bits_rdata_0),
    .io_icache_resp_bits_rdata_1(fe_io_icache_resp_bits_rdata_1),
    .io_icache_resp_bits_respn(fe_io_icache_resp_bits_respn),
    .cache_stall_0(fe_cache_stall_0)
  );
  Backend be ( // @[Core.scala 98:18]
    .clock(be_clock),
    .reset(be_reset),
    .io_fb_bmfs_redirect_kill(be_io_fb_bmfs_redirect_kill),
    .io_fb_bmfs_redirect_pc(be_io_fb_bmfs_redirect_pc),
    .io_fb_bmfs_bpu_v(be_io_fb_bmfs_bpu_v),
    .io_fb_bmfs_bpu_errpr(be_io_fb_bmfs_bpu_errpr),
    .io_fb_bmfs_bpu_pc_br(be_io_fb_bmfs_bpu_pc_br),
    .io_fb_bmfs_bpu_target(be_io_fb_bmfs_bpu_target),
    .io_fb_bmfs_bpu_taken(be_io_fb_bmfs_bpu_taken),
    .io_fb_fmbs_instn(be_io_fb_fmbs_instn),
    .io_fb_fmbs_inst_ops_0(be_io_fb_fmbs_inst_ops_0),
    .io_fb_fmbs_inst_ops_1(be_io_fb_fmbs_inst_ops_1),
    .io_fb_fmbs_please_wait(be_io_fb_fmbs_please_wait),
    .io_dcache_req_valid(be_io_dcache_req_valid),
    .io_dcache_req_bits_addr(be_io_dcache_req_bits_addr),
    .io_dcache_req_bits_wdata(be_io_dcache_req_bits_wdata),
    .io_dcache_req_bits_wen(be_io_dcache_req_bits_wen),
    .io_dcache_req_bits_mtype(be_io_dcache_req_bits_mtype),
    .io_dcache_resp_valid(be_io_dcache_resp_valid),
    .io_dcache_resp_bits_rdata_0(be_io_dcache_resp_bits_rdata_0),
    .io_dcache_resp_bits_rdata_1(be_io_dcache_resp_bits_rdata_1),
    .csrs_mstatus(be_csrs_mstatus),
    .csrs_sstatus(be_csrs_sstatus),
    .csrs_mepc(be_csrs_mepc),
    .csrs_sepc(be_csrs_sepc),
    .csrs_mtval(be_csrs_mtval),
    .csrs_stval(be_csrs_stval),
    .csrs_mtvec(be_csrs_mtvec),
    .csrs_stvec(be_csrs_stvec),
    .csrs_mcause(be_csrs_mcause),
    .csrs_scause(be_csrs_scause),
    .csrs_satp(be_csrs_satp),
    .csrs_mip(be_csrs_mip),
    .csrs_mie(be_csrs_mie),
    .csrs_mscratch(be_csrs_mscratch),
    .csrs_sscratch(be_csrs_sscratch),
    .csrs_mideleg(be_csrs_mideleg),
    .csrs_medeleg(be_csrs_medeleg),
    .istall_0(be_istall_0),
    ._WIRE_4_0_0(be__WIRE_4_0_0),
    ._WIRE_4_0_1(be__WIRE_4_0_1),
    ._WIRE_4_0_2(be__WIRE_4_0_2),
    ._WIRE_1_0_0(be__WIRE_1_0_0),
    ._WIRE_1_0_1(be__WIRE_1_0_1),
    ._WIRE_1_0_2(be__WIRE_1_0_2),
    .difftest_saddr(be_difftest_saddr),
    .current_mode(be_current_mode),
    ._WIRE_0_0(be__WIRE_0_0),
    ._WIRE_0_1(be__WIRE_0_1),
    ._WIRE_0_2(be__WIRE_0_2),
    ._WIRE_0_3(be__WIRE_0_3),
    ._WIRE_0_4(be__WIRE_0_4),
    ._WIRE_0_5(be__WIRE_0_5),
    ._WIRE_0_6(be__WIRE_0_6),
    ._WIRE_0_7(be__WIRE_0_7),
    ._WIRE_0_8(be__WIRE_0_8),
    ._WIRE_0_9(be__WIRE_0_9),
    ._WIRE_0_10(be__WIRE_0_10),
    ._WIRE_0_11(be__WIRE_0_11),
    ._WIRE_0_12(be__WIRE_0_12),
    ._WIRE_0_13(be__WIRE_0_13),
    ._WIRE_0_14(be__WIRE_0_14),
    ._WIRE_0_15(be__WIRE_0_15),
    ._WIRE_0_16(be__WIRE_0_16),
    ._WIRE_0_17(be__WIRE_0_17),
    ._WIRE_0_18(be__WIRE_0_18),
    ._WIRE_0_19(be__WIRE_0_19),
    ._WIRE_0_20(be__WIRE_0_20),
    ._WIRE_0_21(be__WIRE_0_21),
    ._WIRE_0_22(be__WIRE_0_22),
    ._WIRE_0_23(be__WIRE_0_23),
    ._WIRE_0_24(be__WIRE_0_24),
    ._WIRE_0_25(be__WIRE_0_25),
    ._WIRE_0_26(be__WIRE_0_26),
    ._WIRE_0_27(be__WIRE_0_27),
    ._WIRE_0_28(be__WIRE_0_28),
    ._WIRE_0_29(be__WIRE_0_29),
    ._WIRE_0_30(be__WIRE_0_30),
    ._WIRE_0_31(be__WIRE_0_31),
    .dstall_0(be_dstall_0),
    ._WIRE_6_0(be__WIRE_6_0),
    ._WIRE_6_1(be__WIRE_6_1),
    ._WIRE_6_2(be__WIRE_6_2),
    .counter_0(be_counter_0),
    .icache_stall(be_icache_stall),
    .difftest_sval(be_difftest_sval),
    .mduStall_0(be_mduStall_0),
    ._WIRE_3_0_0(be__WIRE_3_0_0),
    ._WIRE_3_0_1(be__WIRE_3_0_1),
    ._WIRE_3_0_2(be__WIRE_3_0_2),
    .common_0(be_common_0),
    ._WIRE_5_0_0(be__WIRE_5_0_0),
    ._WIRE_5_0_1(be__WIRE_5_0_1),
    ._WIRE_5_0_2(be__WIRE_5_0_2),
    .instret_0(be_instret_0),
    ._WIRE_2_0_0(be__WIRE_2_0_0),
    ._WIRE_2_0_1(be__WIRE_2_0_1),
    ._WIRE_2_0_2(be__WIRE_2_0_2),
    .REG_0(be_REG_0),
    .difftest_sync(be_difftest_sync),
    .wbInsts_0_ysyx_debug(be_wbInsts_0_ysyx_debug)
  );
  assign io_icache_req_bits_addr = fe_io_icache_req_bits_addr; // @[Core.scala 103:13]
  assign io_icache_req_bits_mtype = fe_io_icache_req_bits_mtype; // @[Core.scala 103:13]
  assign io_dcache_req_valid = be_io_dcache_req_valid; // @[Core.scala 104:13]
  assign io_dcache_req_bits_addr = be_io_dcache_req_bits_addr; // @[Core.scala 104:13]
  assign io_dcache_req_bits_wdata = be_io_dcache_req_bits_wdata; // @[Core.scala 104:13]
  assign io_dcache_req_bits_wen = be_io_dcache_req_bits_wen; // @[Core.scala 104:13]
  assign io_dcache_req_bits_mtype = be_io_dcache_req_bits_mtype; // @[Core.scala 104:13]
  assign csrs_mstatus = be_csrs_mstatus;
  assign csrs_sstatus = be_csrs_sstatus;
  assign csrs_mepc = be_csrs_mepc;
  assign csrs_sepc = be_csrs_sepc;
  assign csrs_mtval = be_csrs_mtval;
  assign csrs_stval = be_csrs_stval;
  assign csrs_mtvec = be_csrs_mtvec;
  assign csrs_stvec = be_csrs_stvec;
  assign csrs_mcause = be_csrs_mcause;
  assign csrs_scause = be_csrs_scause;
  assign csrs_satp = be_csrs_satp;
  assign csrs_mip = be_csrs_mip;
  assign csrs_mie = be_csrs_mie;
  assign csrs_mscratch = be_csrs_mscratch;
  assign csrs_sscratch = be_csrs_sscratch;
  assign csrs_mideleg = be_csrs_mideleg;
  assign csrs_medeleg = be_csrs_medeleg;
  assign istall = be_istall_0;
  assign _WIRE_4_0 = be__WIRE_4_0_0;
  assign _WIRE_4_1 = be__WIRE_4_0_1;
  assign _WIRE_4_2 = be__WIRE_4_0_2;
  assign _WIRE_1_0 = be__WIRE_1_0_0;
  assign _WIRE_1_1 = be__WIRE_1_0_1;
  assign _WIRE_1_2 = be__WIRE_1_0_2;
  assign current_mode = be_current_mode;
  assign _WIRE__0 = be__WIRE_0_0;
  assign _WIRE__1 = be__WIRE_0_1;
  assign _WIRE__2 = be__WIRE_0_2;
  assign _WIRE__3 = be__WIRE_0_3;
  assign _WIRE__4 = be__WIRE_0_4;
  assign _WIRE__5 = be__WIRE_0_5;
  assign _WIRE__6 = be__WIRE_0_6;
  assign _WIRE__7 = be__WIRE_0_7;
  assign _WIRE__8 = be__WIRE_0_8;
  assign _WIRE__9 = be__WIRE_0_9;
  assign _WIRE__10 = be__WIRE_0_10;
  assign _WIRE__11 = be__WIRE_0_11;
  assign _WIRE__12 = be__WIRE_0_12;
  assign _WIRE__13 = be__WIRE_0_13;
  assign _WIRE__14 = be__WIRE_0_14;
  assign _WIRE__15 = be__WIRE_0_15;
  assign _WIRE__16 = be__WIRE_0_16;
  assign _WIRE__17 = be__WIRE_0_17;
  assign _WIRE__18 = be__WIRE_0_18;
  assign _WIRE__19 = be__WIRE_0_19;
  assign _WIRE__20 = be__WIRE_0_20;
  assign _WIRE__21 = be__WIRE_0_21;
  assign _WIRE__22 = be__WIRE_0_22;
  assign _WIRE__23 = be__WIRE_0_23;
  assign _WIRE__24 = be__WIRE_0_24;
  assign _WIRE__25 = be__WIRE_0_25;
  assign _WIRE__26 = be__WIRE_0_26;
  assign _WIRE__27 = be__WIRE_0_27;
  assign _WIRE__28 = be__WIRE_0_28;
  assign _WIRE__29 = be__WIRE_0_29;
  assign _WIRE__30 = be__WIRE_0_30;
  assign _WIRE__31 = be__WIRE_0_31;
  assign dstall = be_dstall_0;
  assign _WIRE_0_0 = be__WIRE_6_0;
  assign _WIRE_0_1 = be__WIRE_6_1;
  assign _WIRE_0_2 = be__WIRE_6_2;
  assign counter = be_counter_0;
  assign mduStall = be_mduStall_0;
  assign _WIRE_3_0 = be__WIRE_3_0_0;
  assign _WIRE_3_1 = be__WIRE_3_0_1;
  assign _WIRE_3_2 = be__WIRE_3_0_2;
  assign common = be_common_0;
  assign _WIRE_5_0 = be__WIRE_5_0_0;
  assign _WIRE_5_1 = be__WIRE_5_0_1;
  assign _WIRE_5_2 = be__WIRE_5_0_2;
  assign instret = be_instret_0;
  assign _WIRE_2_0 = be__WIRE_2_0_0;
  assign _WIRE_2_1 = be__WIRE_2_0_1;
  assign _WIRE_2_2 = be__WIRE_2_0_2;
  assign REG_0 = be_REG_0;
  assign wbInsts_0_ysyx_debug = be_wbInsts_0_ysyx_debug;
  assign fe_clock = clock;
  assign fe_reset = reset;
  assign fe_io_fb_bmfs_redirect_kill = be_io_fb_bmfs_redirect_kill; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_redirect_pc = be_io_fb_bmfs_redirect_pc; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_bpu_v = be_io_fb_bmfs_bpu_v; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_bpu_errpr = be_io_fb_bmfs_bpu_errpr; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_bpu_pc_br = be_io_fb_bmfs_bpu_pc_br; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_bpu_target = be_io_fb_bmfs_bpu_target; // @[Core.scala 100:12]
  assign fe_io_fb_bmfs_bpu_taken = be_io_fb_bmfs_bpu_taken; // @[Core.scala 100:12]
  assign fe_io_fb_fmbs_please_wait = be_io_fb_fmbs_please_wait; // @[Core.scala 100:12]
  assign fe_io_icache_resp_valid = io_icache_resp_valid; // @[Core.scala 103:13]
  assign fe_io_icache_resp_bits_rdata_0 = io_icache_resp_bits_rdata_0; // @[Core.scala 103:13]
  assign fe_io_icache_resp_bits_rdata_1 = io_icache_resp_bits_rdata_1; // @[Core.scala 103:13]
  assign fe_io_icache_resp_bits_respn = io_icache_resp_bits_respn; // @[Core.scala 103:13]
  assign be_clock = clock;
  assign be_reset = reset;
  assign be_io_fb_fmbs_instn = fe_io_fb_fmbs_instn; // @[Core.scala 100:12]
  assign be_io_fb_fmbs_inst_ops_0 = fe_io_fb_fmbs_inst_ops_0; // @[Core.scala 100:12]
  assign be_io_fb_fmbs_inst_ops_1 = fe_io_fb_fmbs_inst_ops_1; // @[Core.scala 100:12]
  assign be_io_dcache_resp_valid = io_dcache_resp_valid; // @[Core.scala 104:13]
  assign be_io_dcache_resp_bits_rdata_0 = io_dcache_resp_bits_rdata_0; // @[Core.scala 104:13]
  assign be_io_dcache_resp_bits_rdata_1 = io_dcache_resp_bits_rdata_1; // @[Core.scala 104:13]
  assign be_difftest_saddr = difftest_saddr;
  assign be_icache_stall = fe_cache_stall_0;
  assign be_difftest_sval = difftest_sval;
  assign be_difftest_sync = difftest_sync;
endmodule
module SimSinglePortBRAM(
  input          clock,
  input          reset,
  input          io_we,
  input  [8:0]   io_addr,
  input  [255:0] io_din,
  output [255:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [255:0] _RAND_2;
  reg [255:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [255:0] _RAND_5;
  reg [255:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [255:0] _RAND_9;
  reg [255:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [255:0] _RAND_12;
  reg [255:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [255:0] _RAND_16;
  reg [255:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [255:0] _RAND_22;
  reg [255:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [255:0] _RAND_26;
  reg [255:0] _RAND_27;
  reg [255:0] _RAND_28;
  reg [255:0] _RAND_29;
  reg [255:0] _RAND_30;
  reg [255:0] _RAND_31;
  reg [255:0] _RAND_32;
  reg [255:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [255:0] _RAND_35;
  reg [255:0] _RAND_36;
  reg [255:0] _RAND_37;
  reg [255:0] _RAND_38;
  reg [255:0] _RAND_39;
  reg [255:0] _RAND_40;
  reg [255:0] _RAND_41;
  reg [255:0] _RAND_42;
  reg [255:0] _RAND_43;
  reg [255:0] _RAND_44;
  reg [255:0] _RAND_45;
  reg [255:0] _RAND_46;
  reg [255:0] _RAND_47;
  reg [255:0] _RAND_48;
  reg [255:0] _RAND_49;
  reg [255:0] _RAND_50;
  reg [255:0] _RAND_51;
  reg [255:0] _RAND_52;
  reg [255:0] _RAND_53;
  reg [255:0] _RAND_54;
  reg [255:0] _RAND_55;
  reg [255:0] _RAND_56;
  reg [255:0] _RAND_57;
  reg [255:0] _RAND_58;
  reg [255:0] _RAND_59;
  reg [255:0] _RAND_60;
  reg [255:0] _RAND_61;
  reg [255:0] _RAND_62;
  reg [255:0] _RAND_63;
  reg [255:0] _RAND_64;
  reg [255:0] _RAND_65;
  reg [255:0] _RAND_66;
  reg [255:0] _RAND_67;
  reg [255:0] _RAND_68;
  reg [255:0] _RAND_69;
  reg [255:0] _RAND_70;
  reg [255:0] _RAND_71;
  reg [255:0] _RAND_72;
  reg [255:0] _RAND_73;
  reg [255:0] _RAND_74;
  reg [255:0] _RAND_75;
  reg [255:0] _RAND_76;
  reg [255:0] _RAND_77;
  reg [255:0] _RAND_78;
  reg [255:0] _RAND_79;
  reg [255:0] _RAND_80;
  reg [255:0] _RAND_81;
  reg [255:0] _RAND_82;
  reg [255:0] _RAND_83;
  reg [255:0] _RAND_84;
  reg [255:0] _RAND_85;
  reg [255:0] _RAND_86;
  reg [255:0] _RAND_87;
  reg [255:0] _RAND_88;
  reg [255:0] _RAND_89;
  reg [255:0] _RAND_90;
  reg [255:0] _RAND_91;
  reg [255:0] _RAND_92;
  reg [255:0] _RAND_93;
  reg [255:0] _RAND_94;
  reg [255:0] _RAND_95;
  reg [255:0] _RAND_96;
  reg [255:0] _RAND_97;
  reg [255:0] _RAND_98;
  reg [255:0] _RAND_99;
  reg [255:0] _RAND_100;
  reg [255:0] _RAND_101;
  reg [255:0] _RAND_102;
  reg [255:0] _RAND_103;
  reg [255:0] _RAND_104;
  reg [255:0] _RAND_105;
  reg [255:0] _RAND_106;
  reg [255:0] _RAND_107;
  reg [255:0] _RAND_108;
  reg [255:0] _RAND_109;
  reg [255:0] _RAND_110;
  reg [255:0] _RAND_111;
  reg [255:0] _RAND_112;
  reg [255:0] _RAND_113;
  reg [255:0] _RAND_114;
  reg [255:0] _RAND_115;
  reg [255:0] _RAND_116;
  reg [255:0] _RAND_117;
  reg [255:0] _RAND_118;
  reg [255:0] _RAND_119;
  reg [255:0] _RAND_120;
  reg [255:0] _RAND_121;
  reg [255:0] _RAND_122;
  reg [255:0] _RAND_123;
  reg [255:0] _RAND_124;
  reg [255:0] _RAND_125;
  reg [255:0] _RAND_126;
  reg [255:0] _RAND_127;
  reg [255:0] _RAND_128;
  reg [255:0] _RAND_129;
  reg [255:0] _RAND_130;
  reg [255:0] _RAND_131;
  reg [255:0] _RAND_132;
  reg [255:0] _RAND_133;
  reg [255:0] _RAND_134;
  reg [255:0] _RAND_135;
  reg [255:0] _RAND_136;
  reg [255:0] _RAND_137;
  reg [255:0] _RAND_138;
  reg [255:0] _RAND_139;
  reg [255:0] _RAND_140;
  reg [255:0] _RAND_141;
  reg [255:0] _RAND_142;
  reg [255:0] _RAND_143;
  reg [255:0] _RAND_144;
  reg [255:0] _RAND_145;
  reg [255:0] _RAND_146;
  reg [255:0] _RAND_147;
  reg [255:0] _RAND_148;
  reg [255:0] _RAND_149;
  reg [255:0] _RAND_150;
  reg [255:0] _RAND_151;
  reg [255:0] _RAND_152;
  reg [255:0] _RAND_153;
  reg [255:0] _RAND_154;
  reg [255:0] _RAND_155;
  reg [255:0] _RAND_156;
  reg [255:0] _RAND_157;
  reg [255:0] _RAND_158;
  reg [255:0] _RAND_159;
  reg [255:0] _RAND_160;
  reg [255:0] _RAND_161;
  reg [255:0] _RAND_162;
  reg [255:0] _RAND_163;
  reg [255:0] _RAND_164;
  reg [255:0] _RAND_165;
  reg [255:0] _RAND_166;
  reg [255:0] _RAND_167;
  reg [255:0] _RAND_168;
  reg [255:0] _RAND_169;
  reg [255:0] _RAND_170;
  reg [255:0] _RAND_171;
  reg [255:0] _RAND_172;
  reg [255:0] _RAND_173;
  reg [255:0] _RAND_174;
  reg [255:0] _RAND_175;
  reg [255:0] _RAND_176;
  reg [255:0] _RAND_177;
  reg [255:0] _RAND_178;
  reg [255:0] _RAND_179;
  reg [255:0] _RAND_180;
  reg [255:0] _RAND_181;
  reg [255:0] _RAND_182;
  reg [255:0] _RAND_183;
  reg [255:0] _RAND_184;
  reg [255:0] _RAND_185;
  reg [255:0] _RAND_186;
  reg [255:0] _RAND_187;
  reg [255:0] _RAND_188;
  reg [255:0] _RAND_189;
  reg [255:0] _RAND_190;
  reg [255:0] _RAND_191;
  reg [255:0] _RAND_192;
  reg [255:0] _RAND_193;
  reg [255:0] _RAND_194;
  reg [255:0] _RAND_195;
  reg [255:0] _RAND_196;
  reg [255:0] _RAND_197;
  reg [255:0] _RAND_198;
  reg [255:0] _RAND_199;
  reg [255:0] _RAND_200;
  reg [255:0] _RAND_201;
  reg [255:0] _RAND_202;
  reg [255:0] _RAND_203;
  reg [255:0] _RAND_204;
  reg [255:0] _RAND_205;
  reg [255:0] _RAND_206;
  reg [255:0] _RAND_207;
  reg [255:0] _RAND_208;
  reg [255:0] _RAND_209;
  reg [255:0] _RAND_210;
  reg [255:0] _RAND_211;
  reg [255:0] _RAND_212;
  reg [255:0] _RAND_213;
  reg [255:0] _RAND_214;
  reg [255:0] _RAND_215;
  reg [255:0] _RAND_216;
  reg [255:0] _RAND_217;
  reg [255:0] _RAND_218;
  reg [255:0] _RAND_219;
  reg [255:0] _RAND_220;
  reg [255:0] _RAND_221;
  reg [255:0] _RAND_222;
  reg [255:0] _RAND_223;
  reg [255:0] _RAND_224;
  reg [255:0] _RAND_225;
  reg [255:0] _RAND_226;
  reg [255:0] _RAND_227;
  reg [255:0] _RAND_228;
  reg [255:0] _RAND_229;
  reg [255:0] _RAND_230;
  reg [255:0] _RAND_231;
  reg [255:0] _RAND_232;
  reg [255:0] _RAND_233;
  reg [255:0] _RAND_234;
  reg [255:0] _RAND_235;
  reg [255:0] _RAND_236;
  reg [255:0] _RAND_237;
  reg [255:0] _RAND_238;
  reg [255:0] _RAND_239;
  reg [255:0] _RAND_240;
  reg [255:0] _RAND_241;
  reg [255:0] _RAND_242;
  reg [255:0] _RAND_243;
  reg [255:0] _RAND_244;
  reg [255:0] _RAND_245;
  reg [255:0] _RAND_246;
  reg [255:0] _RAND_247;
  reg [255:0] _RAND_248;
  reg [255:0] _RAND_249;
  reg [255:0] _RAND_250;
  reg [255:0] _RAND_251;
  reg [255:0] _RAND_252;
  reg [255:0] _RAND_253;
  reg [255:0] _RAND_254;
  reg [255:0] _RAND_255;
  reg [255:0] _RAND_256;
  reg [255:0] _RAND_257;
  reg [255:0] _RAND_258;
  reg [255:0] _RAND_259;
  reg [255:0] _RAND_260;
  reg [255:0] _RAND_261;
  reg [255:0] _RAND_262;
  reg [255:0] _RAND_263;
  reg [255:0] _RAND_264;
  reg [255:0] _RAND_265;
  reg [255:0] _RAND_266;
  reg [255:0] _RAND_267;
  reg [255:0] _RAND_268;
  reg [255:0] _RAND_269;
  reg [255:0] _RAND_270;
  reg [255:0] _RAND_271;
  reg [255:0] _RAND_272;
  reg [255:0] _RAND_273;
  reg [255:0] _RAND_274;
  reg [255:0] _RAND_275;
  reg [255:0] _RAND_276;
  reg [255:0] _RAND_277;
  reg [255:0] _RAND_278;
  reg [255:0] _RAND_279;
  reg [255:0] _RAND_280;
  reg [255:0] _RAND_281;
  reg [255:0] _RAND_282;
  reg [255:0] _RAND_283;
  reg [255:0] _RAND_284;
  reg [255:0] _RAND_285;
  reg [255:0] _RAND_286;
  reg [255:0] _RAND_287;
  reg [255:0] _RAND_288;
  reg [255:0] _RAND_289;
  reg [255:0] _RAND_290;
  reg [255:0] _RAND_291;
  reg [255:0] _RAND_292;
  reg [255:0] _RAND_293;
  reg [255:0] _RAND_294;
  reg [255:0] _RAND_295;
  reg [255:0] _RAND_296;
  reg [255:0] _RAND_297;
  reg [255:0] _RAND_298;
  reg [255:0] _RAND_299;
  reg [255:0] _RAND_300;
  reg [255:0] _RAND_301;
  reg [255:0] _RAND_302;
  reg [255:0] _RAND_303;
  reg [255:0] _RAND_304;
  reg [255:0] _RAND_305;
  reg [255:0] _RAND_306;
  reg [255:0] _RAND_307;
  reg [255:0] _RAND_308;
  reg [255:0] _RAND_309;
  reg [255:0] _RAND_310;
  reg [255:0] _RAND_311;
  reg [255:0] _RAND_312;
  reg [255:0] _RAND_313;
  reg [255:0] _RAND_314;
  reg [255:0] _RAND_315;
  reg [255:0] _RAND_316;
  reg [255:0] _RAND_317;
  reg [255:0] _RAND_318;
  reg [255:0] _RAND_319;
  reg [255:0] _RAND_320;
  reg [255:0] _RAND_321;
  reg [255:0] _RAND_322;
  reg [255:0] _RAND_323;
  reg [255:0] _RAND_324;
  reg [255:0] _RAND_325;
  reg [255:0] _RAND_326;
  reg [255:0] _RAND_327;
  reg [255:0] _RAND_328;
  reg [255:0] _RAND_329;
  reg [255:0] _RAND_330;
  reg [255:0] _RAND_331;
  reg [255:0] _RAND_332;
  reg [255:0] _RAND_333;
  reg [255:0] _RAND_334;
  reg [255:0] _RAND_335;
  reg [255:0] _RAND_336;
  reg [255:0] _RAND_337;
  reg [255:0] _RAND_338;
  reg [255:0] _RAND_339;
  reg [255:0] _RAND_340;
  reg [255:0] _RAND_341;
  reg [255:0] _RAND_342;
  reg [255:0] _RAND_343;
  reg [255:0] _RAND_344;
  reg [255:0] _RAND_345;
  reg [255:0] _RAND_346;
  reg [255:0] _RAND_347;
  reg [255:0] _RAND_348;
  reg [255:0] _RAND_349;
  reg [255:0] _RAND_350;
  reg [255:0] _RAND_351;
  reg [255:0] _RAND_352;
  reg [255:0] _RAND_353;
  reg [255:0] _RAND_354;
  reg [255:0] _RAND_355;
  reg [255:0] _RAND_356;
  reg [255:0] _RAND_357;
  reg [255:0] _RAND_358;
  reg [255:0] _RAND_359;
  reg [255:0] _RAND_360;
  reg [255:0] _RAND_361;
  reg [255:0] _RAND_362;
  reg [255:0] _RAND_363;
  reg [255:0] _RAND_364;
  reg [255:0] _RAND_365;
  reg [255:0] _RAND_366;
  reg [255:0] _RAND_367;
  reg [255:0] _RAND_368;
  reg [255:0] _RAND_369;
  reg [255:0] _RAND_370;
  reg [255:0] _RAND_371;
  reg [255:0] _RAND_372;
  reg [255:0] _RAND_373;
  reg [255:0] _RAND_374;
  reg [255:0] _RAND_375;
  reg [255:0] _RAND_376;
  reg [255:0] _RAND_377;
  reg [255:0] _RAND_378;
  reg [255:0] _RAND_379;
  reg [255:0] _RAND_380;
  reg [255:0] _RAND_381;
  reg [255:0] _RAND_382;
  reg [255:0] _RAND_383;
  reg [255:0] _RAND_384;
  reg [255:0] _RAND_385;
  reg [255:0] _RAND_386;
  reg [255:0] _RAND_387;
  reg [255:0] _RAND_388;
  reg [255:0] _RAND_389;
  reg [255:0] _RAND_390;
  reg [255:0] _RAND_391;
  reg [255:0] _RAND_392;
  reg [255:0] _RAND_393;
  reg [255:0] _RAND_394;
  reg [255:0] _RAND_395;
  reg [255:0] _RAND_396;
  reg [255:0] _RAND_397;
  reg [255:0] _RAND_398;
  reg [255:0] _RAND_399;
  reg [255:0] _RAND_400;
  reg [255:0] _RAND_401;
  reg [255:0] _RAND_402;
  reg [255:0] _RAND_403;
  reg [255:0] _RAND_404;
  reg [255:0] _RAND_405;
  reg [255:0] _RAND_406;
  reg [255:0] _RAND_407;
  reg [255:0] _RAND_408;
  reg [255:0] _RAND_409;
  reg [255:0] _RAND_410;
  reg [255:0] _RAND_411;
  reg [255:0] _RAND_412;
  reg [255:0] _RAND_413;
  reg [255:0] _RAND_414;
  reg [255:0] _RAND_415;
  reg [255:0] _RAND_416;
  reg [255:0] _RAND_417;
  reg [255:0] _RAND_418;
  reg [255:0] _RAND_419;
  reg [255:0] _RAND_420;
  reg [255:0] _RAND_421;
  reg [255:0] _RAND_422;
  reg [255:0] _RAND_423;
  reg [255:0] _RAND_424;
  reg [255:0] _RAND_425;
  reg [255:0] _RAND_426;
  reg [255:0] _RAND_427;
  reg [255:0] _RAND_428;
  reg [255:0] _RAND_429;
  reg [255:0] _RAND_430;
  reg [255:0] _RAND_431;
  reg [255:0] _RAND_432;
  reg [255:0] _RAND_433;
  reg [255:0] _RAND_434;
  reg [255:0] _RAND_435;
  reg [255:0] _RAND_436;
  reg [255:0] _RAND_437;
  reg [255:0] _RAND_438;
  reg [255:0] _RAND_439;
  reg [255:0] _RAND_440;
  reg [255:0] _RAND_441;
  reg [255:0] _RAND_442;
  reg [255:0] _RAND_443;
  reg [255:0] _RAND_444;
  reg [255:0] _RAND_445;
  reg [255:0] _RAND_446;
  reg [255:0] _RAND_447;
  reg [255:0] _RAND_448;
  reg [255:0] _RAND_449;
  reg [255:0] _RAND_450;
  reg [255:0] _RAND_451;
  reg [255:0] _RAND_452;
  reg [255:0] _RAND_453;
  reg [255:0] _RAND_454;
  reg [255:0] _RAND_455;
  reg [255:0] _RAND_456;
  reg [255:0] _RAND_457;
  reg [255:0] _RAND_458;
  reg [255:0] _RAND_459;
  reg [255:0] _RAND_460;
  reg [255:0] _RAND_461;
  reg [255:0] _RAND_462;
  reg [255:0] _RAND_463;
  reg [255:0] _RAND_464;
  reg [255:0] _RAND_465;
  reg [255:0] _RAND_466;
  reg [255:0] _RAND_467;
  reg [255:0] _RAND_468;
  reg [255:0] _RAND_469;
  reg [255:0] _RAND_470;
  reg [255:0] _RAND_471;
  reg [255:0] _RAND_472;
  reg [255:0] _RAND_473;
  reg [255:0] _RAND_474;
  reg [255:0] _RAND_475;
  reg [255:0] _RAND_476;
  reg [255:0] _RAND_477;
  reg [255:0] _RAND_478;
  reg [255:0] _RAND_479;
  reg [255:0] _RAND_480;
  reg [255:0] _RAND_481;
  reg [255:0] _RAND_482;
  reg [255:0] _RAND_483;
  reg [255:0] _RAND_484;
  reg [255:0] _RAND_485;
  reg [255:0] _RAND_486;
  reg [255:0] _RAND_487;
  reg [255:0] _RAND_488;
  reg [255:0] _RAND_489;
  reg [255:0] _RAND_490;
  reg [255:0] _RAND_491;
  reg [255:0] _RAND_492;
  reg [255:0] _RAND_493;
  reg [255:0] _RAND_494;
  reg [255:0] _RAND_495;
  reg [255:0] _RAND_496;
  reg [255:0] _RAND_497;
  reg [255:0] _RAND_498;
  reg [255:0] _RAND_499;
  reg [255:0] _RAND_500;
  reg [255:0] _RAND_501;
  reg [255:0] _RAND_502;
  reg [255:0] _RAND_503;
  reg [255:0] _RAND_504;
  reg [255:0] _RAND_505;
  reg [255:0] _RAND_506;
  reg [255:0] _RAND_507;
  reg [255:0] _RAND_508;
  reg [255:0] _RAND_509;
  reg [255:0] _RAND_510;
  reg [255:0] _RAND_511;
  reg [255:0] _RAND_512;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] mem_0; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_1; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_2; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_3; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_4; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_5; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_6; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_7; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_8; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_9; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_10; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_11; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_12; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_13; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_14; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_15; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_16; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_17; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_18; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_19; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_20; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_21; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_22; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_23; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_24; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_25; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_26; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_27; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_28; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_29; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_30; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_31; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_32; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_33; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_34; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_35; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_36; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_37; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_38; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_39; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_40; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_41; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_42; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_43; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_44; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_45; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_46; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_47; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_48; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_49; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_50; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_51; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_52; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_53; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_54; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_55; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_56; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_57; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_58; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_59; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_60; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_61; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_62; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_63; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_64; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_65; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_66; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_67; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_68; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_69; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_70; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_71; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_72; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_73; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_74; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_75; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_76; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_77; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_78; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_79; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_80; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_81; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_82; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_83; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_84; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_85; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_86; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_87; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_88; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_89; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_90; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_91; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_92; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_93; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_94; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_95; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_96; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_97; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_98; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_99; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_100; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_101; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_102; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_103; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_104; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_105; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_106; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_107; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_108; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_109; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_110; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_111; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_112; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_113; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_114; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_115; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_116; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_117; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_118; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_119; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_120; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_121; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_122; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_123; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_124; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_125; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_126; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_127; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_128; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_129; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_130; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_131; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_132; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_133; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_134; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_135; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_136; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_137; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_138; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_139; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_140; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_141; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_142; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_143; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_144; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_145; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_146; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_147; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_148; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_149; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_150; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_151; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_152; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_153; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_154; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_155; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_156; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_157; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_158; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_159; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_160; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_161; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_162; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_163; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_164; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_165; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_166; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_167; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_168; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_169; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_170; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_171; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_172; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_173; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_174; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_175; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_176; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_177; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_178; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_179; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_180; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_181; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_182; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_183; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_184; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_185; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_186; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_187; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_188; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_189; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_190; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_191; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_192; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_193; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_194; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_195; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_196; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_197; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_198; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_199; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_200; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_201; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_202; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_203; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_204; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_205; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_206; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_207; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_208; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_209; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_210; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_211; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_212; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_213; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_214; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_215; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_216; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_217; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_218; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_219; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_220; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_221; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_222; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_223; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_224; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_225; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_226; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_227; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_228; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_229; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_230; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_231; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_232; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_233; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_234; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_235; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_236; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_237; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_238; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_239; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_240; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_241; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_242; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_243; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_244; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_245; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_246; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_247; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_248; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_249; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_250; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_251; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_252; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_253; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_254; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_255; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_256; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_257; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_258; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_259; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_260; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_261; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_262; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_263; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_264; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_265; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_266; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_267; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_268; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_269; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_270; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_271; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_272; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_273; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_274; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_275; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_276; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_277; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_278; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_279; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_280; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_281; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_282; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_283; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_284; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_285; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_286; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_287; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_288; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_289; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_290; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_291; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_292; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_293; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_294; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_295; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_296; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_297; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_298; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_299; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_300; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_301; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_302; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_303; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_304; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_305; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_306; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_307; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_308; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_309; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_310; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_311; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_312; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_313; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_314; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_315; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_316; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_317; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_318; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_319; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_320; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_321; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_322; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_323; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_324; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_325; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_326; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_327; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_328; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_329; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_330; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_331; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_332; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_333; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_334; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_335; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_336; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_337; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_338; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_339; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_340; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_341; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_342; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_343; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_344; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_345; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_346; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_347; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_348; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_349; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_350; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_351; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_352; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_353; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_354; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_355; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_356; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_357; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_358; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_359; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_360; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_361; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_362; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_363; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_364; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_365; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_366; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_367; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_368; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_369; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_370; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_371; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_372; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_373; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_374; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_375; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_376; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_377; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_378; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_379; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_380; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_381; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_382; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_383; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_384; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_385; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_386; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_387; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_388; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_389; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_390; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_391; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_392; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_393; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_394; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_395; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_396; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_397; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_398; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_399; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_400; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_401; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_402; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_403; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_404; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_405; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_406; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_407; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_408; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_409; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_410; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_411; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_412; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_413; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_414; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_415; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_416; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_417; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_418; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_419; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_420; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_421; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_422; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_423; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_424; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_425; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_426; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_427; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_428; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_429; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_430; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_431; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_432; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_433; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_434; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_435; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_436; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_437; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_438; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_439; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_440; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_441; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_442; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_443; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_444; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_445; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_446; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_447; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_448; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_449; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_450; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_451; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_452; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_453; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_454; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_455; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_456; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_457; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_458; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_459; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_460; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_461; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_462; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_463; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_464; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_465; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_466; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_467; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_468; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_469; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_470; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_471; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_472; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_473; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_474; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_475; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_476; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_477; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_478; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_479; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_480; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_481; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_482; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_483; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_484; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_485; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_486; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_487; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_488; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_489; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_490; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_491; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_492; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_493; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_494; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_495; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_496; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_497; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_498; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_499; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_500; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_501; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_502; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_503; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_504; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_505; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_506; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_507; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_508; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_509; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_510; // @[RAMWrapper.scala 286:20]
  reg [255:0] mem_511; // @[RAMWrapper.scala 286:20]
  reg [255:0] io_dout_REG; // @[RAMWrapper.scala 288:21]
  wire [255:0] _GEN_1 = 9'h1 == io_addr ? mem_1 : mem_0; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_2 = 9'h2 == io_addr ? mem_2 : _GEN_1; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_3 = 9'h3 == io_addr ? mem_3 : _GEN_2; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_4 = 9'h4 == io_addr ? mem_4 : _GEN_3; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_5 = 9'h5 == io_addr ? mem_5 : _GEN_4; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_6 = 9'h6 == io_addr ? mem_6 : _GEN_5; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_7 = 9'h7 == io_addr ? mem_7 : _GEN_6; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_8 = 9'h8 == io_addr ? mem_8 : _GEN_7; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_9 = 9'h9 == io_addr ? mem_9 : _GEN_8; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_10 = 9'ha == io_addr ? mem_10 : _GEN_9; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_11 = 9'hb == io_addr ? mem_11 : _GEN_10; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_12 = 9'hc == io_addr ? mem_12 : _GEN_11; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_13 = 9'hd == io_addr ? mem_13 : _GEN_12; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_14 = 9'he == io_addr ? mem_14 : _GEN_13; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_15 = 9'hf == io_addr ? mem_15 : _GEN_14; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_16 = 9'h10 == io_addr ? mem_16 : _GEN_15; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_17 = 9'h11 == io_addr ? mem_17 : _GEN_16; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_18 = 9'h12 == io_addr ? mem_18 : _GEN_17; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_19 = 9'h13 == io_addr ? mem_19 : _GEN_18; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_20 = 9'h14 == io_addr ? mem_20 : _GEN_19; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_21 = 9'h15 == io_addr ? mem_21 : _GEN_20; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_22 = 9'h16 == io_addr ? mem_22 : _GEN_21; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_23 = 9'h17 == io_addr ? mem_23 : _GEN_22; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_24 = 9'h18 == io_addr ? mem_24 : _GEN_23; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_25 = 9'h19 == io_addr ? mem_25 : _GEN_24; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_26 = 9'h1a == io_addr ? mem_26 : _GEN_25; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_27 = 9'h1b == io_addr ? mem_27 : _GEN_26; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_28 = 9'h1c == io_addr ? mem_28 : _GEN_27; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_29 = 9'h1d == io_addr ? mem_29 : _GEN_28; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_30 = 9'h1e == io_addr ? mem_30 : _GEN_29; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_31 = 9'h1f == io_addr ? mem_31 : _GEN_30; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_32 = 9'h20 == io_addr ? mem_32 : _GEN_31; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_33 = 9'h21 == io_addr ? mem_33 : _GEN_32; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_34 = 9'h22 == io_addr ? mem_34 : _GEN_33; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_35 = 9'h23 == io_addr ? mem_35 : _GEN_34; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_36 = 9'h24 == io_addr ? mem_36 : _GEN_35; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_37 = 9'h25 == io_addr ? mem_37 : _GEN_36; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_38 = 9'h26 == io_addr ? mem_38 : _GEN_37; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_39 = 9'h27 == io_addr ? mem_39 : _GEN_38; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_40 = 9'h28 == io_addr ? mem_40 : _GEN_39; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_41 = 9'h29 == io_addr ? mem_41 : _GEN_40; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_42 = 9'h2a == io_addr ? mem_42 : _GEN_41; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_43 = 9'h2b == io_addr ? mem_43 : _GEN_42; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_44 = 9'h2c == io_addr ? mem_44 : _GEN_43; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_45 = 9'h2d == io_addr ? mem_45 : _GEN_44; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_46 = 9'h2e == io_addr ? mem_46 : _GEN_45; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_47 = 9'h2f == io_addr ? mem_47 : _GEN_46; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_48 = 9'h30 == io_addr ? mem_48 : _GEN_47; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_49 = 9'h31 == io_addr ? mem_49 : _GEN_48; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_50 = 9'h32 == io_addr ? mem_50 : _GEN_49; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_51 = 9'h33 == io_addr ? mem_51 : _GEN_50; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_52 = 9'h34 == io_addr ? mem_52 : _GEN_51; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_53 = 9'h35 == io_addr ? mem_53 : _GEN_52; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_54 = 9'h36 == io_addr ? mem_54 : _GEN_53; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_55 = 9'h37 == io_addr ? mem_55 : _GEN_54; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_56 = 9'h38 == io_addr ? mem_56 : _GEN_55; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_57 = 9'h39 == io_addr ? mem_57 : _GEN_56; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_58 = 9'h3a == io_addr ? mem_58 : _GEN_57; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_59 = 9'h3b == io_addr ? mem_59 : _GEN_58; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_60 = 9'h3c == io_addr ? mem_60 : _GEN_59; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_61 = 9'h3d == io_addr ? mem_61 : _GEN_60; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_62 = 9'h3e == io_addr ? mem_62 : _GEN_61; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_63 = 9'h3f == io_addr ? mem_63 : _GEN_62; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_64 = 9'h40 == io_addr ? mem_64 : _GEN_63; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_65 = 9'h41 == io_addr ? mem_65 : _GEN_64; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_66 = 9'h42 == io_addr ? mem_66 : _GEN_65; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_67 = 9'h43 == io_addr ? mem_67 : _GEN_66; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_68 = 9'h44 == io_addr ? mem_68 : _GEN_67; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_69 = 9'h45 == io_addr ? mem_69 : _GEN_68; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_70 = 9'h46 == io_addr ? mem_70 : _GEN_69; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_71 = 9'h47 == io_addr ? mem_71 : _GEN_70; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_72 = 9'h48 == io_addr ? mem_72 : _GEN_71; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_73 = 9'h49 == io_addr ? mem_73 : _GEN_72; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_74 = 9'h4a == io_addr ? mem_74 : _GEN_73; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_75 = 9'h4b == io_addr ? mem_75 : _GEN_74; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_76 = 9'h4c == io_addr ? mem_76 : _GEN_75; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_77 = 9'h4d == io_addr ? mem_77 : _GEN_76; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_78 = 9'h4e == io_addr ? mem_78 : _GEN_77; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_79 = 9'h4f == io_addr ? mem_79 : _GEN_78; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_80 = 9'h50 == io_addr ? mem_80 : _GEN_79; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_81 = 9'h51 == io_addr ? mem_81 : _GEN_80; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_82 = 9'h52 == io_addr ? mem_82 : _GEN_81; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_83 = 9'h53 == io_addr ? mem_83 : _GEN_82; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_84 = 9'h54 == io_addr ? mem_84 : _GEN_83; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_85 = 9'h55 == io_addr ? mem_85 : _GEN_84; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_86 = 9'h56 == io_addr ? mem_86 : _GEN_85; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_87 = 9'h57 == io_addr ? mem_87 : _GEN_86; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_88 = 9'h58 == io_addr ? mem_88 : _GEN_87; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_89 = 9'h59 == io_addr ? mem_89 : _GEN_88; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_90 = 9'h5a == io_addr ? mem_90 : _GEN_89; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_91 = 9'h5b == io_addr ? mem_91 : _GEN_90; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_92 = 9'h5c == io_addr ? mem_92 : _GEN_91; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_93 = 9'h5d == io_addr ? mem_93 : _GEN_92; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_94 = 9'h5e == io_addr ? mem_94 : _GEN_93; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_95 = 9'h5f == io_addr ? mem_95 : _GEN_94; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_96 = 9'h60 == io_addr ? mem_96 : _GEN_95; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_97 = 9'h61 == io_addr ? mem_97 : _GEN_96; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_98 = 9'h62 == io_addr ? mem_98 : _GEN_97; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_99 = 9'h63 == io_addr ? mem_99 : _GEN_98; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_100 = 9'h64 == io_addr ? mem_100 : _GEN_99; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_101 = 9'h65 == io_addr ? mem_101 : _GEN_100; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_102 = 9'h66 == io_addr ? mem_102 : _GEN_101; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_103 = 9'h67 == io_addr ? mem_103 : _GEN_102; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_104 = 9'h68 == io_addr ? mem_104 : _GEN_103; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_105 = 9'h69 == io_addr ? mem_105 : _GEN_104; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_106 = 9'h6a == io_addr ? mem_106 : _GEN_105; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_107 = 9'h6b == io_addr ? mem_107 : _GEN_106; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_108 = 9'h6c == io_addr ? mem_108 : _GEN_107; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_109 = 9'h6d == io_addr ? mem_109 : _GEN_108; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_110 = 9'h6e == io_addr ? mem_110 : _GEN_109; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_111 = 9'h6f == io_addr ? mem_111 : _GEN_110; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_112 = 9'h70 == io_addr ? mem_112 : _GEN_111; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_113 = 9'h71 == io_addr ? mem_113 : _GEN_112; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_114 = 9'h72 == io_addr ? mem_114 : _GEN_113; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_115 = 9'h73 == io_addr ? mem_115 : _GEN_114; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_116 = 9'h74 == io_addr ? mem_116 : _GEN_115; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_117 = 9'h75 == io_addr ? mem_117 : _GEN_116; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_118 = 9'h76 == io_addr ? mem_118 : _GEN_117; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_119 = 9'h77 == io_addr ? mem_119 : _GEN_118; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_120 = 9'h78 == io_addr ? mem_120 : _GEN_119; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_121 = 9'h79 == io_addr ? mem_121 : _GEN_120; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_122 = 9'h7a == io_addr ? mem_122 : _GEN_121; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_123 = 9'h7b == io_addr ? mem_123 : _GEN_122; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_124 = 9'h7c == io_addr ? mem_124 : _GEN_123; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_125 = 9'h7d == io_addr ? mem_125 : _GEN_124; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_126 = 9'h7e == io_addr ? mem_126 : _GEN_125; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_127 = 9'h7f == io_addr ? mem_127 : _GEN_126; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_128 = 9'h80 == io_addr ? mem_128 : _GEN_127; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_129 = 9'h81 == io_addr ? mem_129 : _GEN_128; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_130 = 9'h82 == io_addr ? mem_130 : _GEN_129; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_131 = 9'h83 == io_addr ? mem_131 : _GEN_130; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_132 = 9'h84 == io_addr ? mem_132 : _GEN_131; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_133 = 9'h85 == io_addr ? mem_133 : _GEN_132; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_134 = 9'h86 == io_addr ? mem_134 : _GEN_133; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_135 = 9'h87 == io_addr ? mem_135 : _GEN_134; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_136 = 9'h88 == io_addr ? mem_136 : _GEN_135; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_137 = 9'h89 == io_addr ? mem_137 : _GEN_136; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_138 = 9'h8a == io_addr ? mem_138 : _GEN_137; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_139 = 9'h8b == io_addr ? mem_139 : _GEN_138; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_140 = 9'h8c == io_addr ? mem_140 : _GEN_139; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_141 = 9'h8d == io_addr ? mem_141 : _GEN_140; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_142 = 9'h8e == io_addr ? mem_142 : _GEN_141; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_143 = 9'h8f == io_addr ? mem_143 : _GEN_142; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_144 = 9'h90 == io_addr ? mem_144 : _GEN_143; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_145 = 9'h91 == io_addr ? mem_145 : _GEN_144; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_146 = 9'h92 == io_addr ? mem_146 : _GEN_145; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_147 = 9'h93 == io_addr ? mem_147 : _GEN_146; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_148 = 9'h94 == io_addr ? mem_148 : _GEN_147; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_149 = 9'h95 == io_addr ? mem_149 : _GEN_148; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_150 = 9'h96 == io_addr ? mem_150 : _GEN_149; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_151 = 9'h97 == io_addr ? mem_151 : _GEN_150; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_152 = 9'h98 == io_addr ? mem_152 : _GEN_151; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_153 = 9'h99 == io_addr ? mem_153 : _GEN_152; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_154 = 9'h9a == io_addr ? mem_154 : _GEN_153; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_155 = 9'h9b == io_addr ? mem_155 : _GEN_154; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_156 = 9'h9c == io_addr ? mem_156 : _GEN_155; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_157 = 9'h9d == io_addr ? mem_157 : _GEN_156; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_158 = 9'h9e == io_addr ? mem_158 : _GEN_157; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_159 = 9'h9f == io_addr ? mem_159 : _GEN_158; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_160 = 9'ha0 == io_addr ? mem_160 : _GEN_159; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_161 = 9'ha1 == io_addr ? mem_161 : _GEN_160; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_162 = 9'ha2 == io_addr ? mem_162 : _GEN_161; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_163 = 9'ha3 == io_addr ? mem_163 : _GEN_162; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_164 = 9'ha4 == io_addr ? mem_164 : _GEN_163; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_165 = 9'ha5 == io_addr ? mem_165 : _GEN_164; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_166 = 9'ha6 == io_addr ? mem_166 : _GEN_165; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_167 = 9'ha7 == io_addr ? mem_167 : _GEN_166; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_168 = 9'ha8 == io_addr ? mem_168 : _GEN_167; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_169 = 9'ha9 == io_addr ? mem_169 : _GEN_168; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_170 = 9'haa == io_addr ? mem_170 : _GEN_169; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_171 = 9'hab == io_addr ? mem_171 : _GEN_170; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_172 = 9'hac == io_addr ? mem_172 : _GEN_171; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_173 = 9'had == io_addr ? mem_173 : _GEN_172; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_174 = 9'hae == io_addr ? mem_174 : _GEN_173; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_175 = 9'haf == io_addr ? mem_175 : _GEN_174; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_176 = 9'hb0 == io_addr ? mem_176 : _GEN_175; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_177 = 9'hb1 == io_addr ? mem_177 : _GEN_176; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_178 = 9'hb2 == io_addr ? mem_178 : _GEN_177; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_179 = 9'hb3 == io_addr ? mem_179 : _GEN_178; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_180 = 9'hb4 == io_addr ? mem_180 : _GEN_179; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_181 = 9'hb5 == io_addr ? mem_181 : _GEN_180; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_182 = 9'hb6 == io_addr ? mem_182 : _GEN_181; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_183 = 9'hb7 == io_addr ? mem_183 : _GEN_182; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_184 = 9'hb8 == io_addr ? mem_184 : _GEN_183; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_185 = 9'hb9 == io_addr ? mem_185 : _GEN_184; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_186 = 9'hba == io_addr ? mem_186 : _GEN_185; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_187 = 9'hbb == io_addr ? mem_187 : _GEN_186; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_188 = 9'hbc == io_addr ? mem_188 : _GEN_187; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_189 = 9'hbd == io_addr ? mem_189 : _GEN_188; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_190 = 9'hbe == io_addr ? mem_190 : _GEN_189; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_191 = 9'hbf == io_addr ? mem_191 : _GEN_190; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_192 = 9'hc0 == io_addr ? mem_192 : _GEN_191; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_193 = 9'hc1 == io_addr ? mem_193 : _GEN_192; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_194 = 9'hc2 == io_addr ? mem_194 : _GEN_193; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_195 = 9'hc3 == io_addr ? mem_195 : _GEN_194; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_196 = 9'hc4 == io_addr ? mem_196 : _GEN_195; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_197 = 9'hc5 == io_addr ? mem_197 : _GEN_196; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_198 = 9'hc6 == io_addr ? mem_198 : _GEN_197; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_199 = 9'hc7 == io_addr ? mem_199 : _GEN_198; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_200 = 9'hc8 == io_addr ? mem_200 : _GEN_199; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_201 = 9'hc9 == io_addr ? mem_201 : _GEN_200; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_202 = 9'hca == io_addr ? mem_202 : _GEN_201; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_203 = 9'hcb == io_addr ? mem_203 : _GEN_202; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_204 = 9'hcc == io_addr ? mem_204 : _GEN_203; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_205 = 9'hcd == io_addr ? mem_205 : _GEN_204; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_206 = 9'hce == io_addr ? mem_206 : _GEN_205; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_207 = 9'hcf == io_addr ? mem_207 : _GEN_206; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_208 = 9'hd0 == io_addr ? mem_208 : _GEN_207; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_209 = 9'hd1 == io_addr ? mem_209 : _GEN_208; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_210 = 9'hd2 == io_addr ? mem_210 : _GEN_209; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_211 = 9'hd3 == io_addr ? mem_211 : _GEN_210; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_212 = 9'hd4 == io_addr ? mem_212 : _GEN_211; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_213 = 9'hd5 == io_addr ? mem_213 : _GEN_212; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_214 = 9'hd6 == io_addr ? mem_214 : _GEN_213; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_215 = 9'hd7 == io_addr ? mem_215 : _GEN_214; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_216 = 9'hd8 == io_addr ? mem_216 : _GEN_215; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_217 = 9'hd9 == io_addr ? mem_217 : _GEN_216; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_218 = 9'hda == io_addr ? mem_218 : _GEN_217; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_219 = 9'hdb == io_addr ? mem_219 : _GEN_218; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_220 = 9'hdc == io_addr ? mem_220 : _GEN_219; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_221 = 9'hdd == io_addr ? mem_221 : _GEN_220; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_222 = 9'hde == io_addr ? mem_222 : _GEN_221; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_223 = 9'hdf == io_addr ? mem_223 : _GEN_222; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_224 = 9'he0 == io_addr ? mem_224 : _GEN_223; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_225 = 9'he1 == io_addr ? mem_225 : _GEN_224; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_226 = 9'he2 == io_addr ? mem_226 : _GEN_225; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_227 = 9'he3 == io_addr ? mem_227 : _GEN_226; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_228 = 9'he4 == io_addr ? mem_228 : _GEN_227; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_229 = 9'he5 == io_addr ? mem_229 : _GEN_228; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_230 = 9'he6 == io_addr ? mem_230 : _GEN_229; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_231 = 9'he7 == io_addr ? mem_231 : _GEN_230; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_232 = 9'he8 == io_addr ? mem_232 : _GEN_231; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_233 = 9'he9 == io_addr ? mem_233 : _GEN_232; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_234 = 9'hea == io_addr ? mem_234 : _GEN_233; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_235 = 9'heb == io_addr ? mem_235 : _GEN_234; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_236 = 9'hec == io_addr ? mem_236 : _GEN_235; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_237 = 9'hed == io_addr ? mem_237 : _GEN_236; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_238 = 9'hee == io_addr ? mem_238 : _GEN_237; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_239 = 9'hef == io_addr ? mem_239 : _GEN_238; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_240 = 9'hf0 == io_addr ? mem_240 : _GEN_239; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_241 = 9'hf1 == io_addr ? mem_241 : _GEN_240; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_242 = 9'hf2 == io_addr ? mem_242 : _GEN_241; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_243 = 9'hf3 == io_addr ? mem_243 : _GEN_242; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_244 = 9'hf4 == io_addr ? mem_244 : _GEN_243; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_245 = 9'hf5 == io_addr ? mem_245 : _GEN_244; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_246 = 9'hf6 == io_addr ? mem_246 : _GEN_245; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_247 = 9'hf7 == io_addr ? mem_247 : _GEN_246; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_248 = 9'hf8 == io_addr ? mem_248 : _GEN_247; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_249 = 9'hf9 == io_addr ? mem_249 : _GEN_248; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_250 = 9'hfa == io_addr ? mem_250 : _GEN_249; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_251 = 9'hfb == io_addr ? mem_251 : _GEN_250; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_252 = 9'hfc == io_addr ? mem_252 : _GEN_251; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_253 = 9'hfd == io_addr ? mem_253 : _GEN_252; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_254 = 9'hfe == io_addr ? mem_254 : _GEN_253; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_255 = 9'hff == io_addr ? mem_255 : _GEN_254; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_256 = 9'h100 == io_addr ? mem_256 : _GEN_255; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_257 = 9'h101 == io_addr ? mem_257 : _GEN_256; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_258 = 9'h102 == io_addr ? mem_258 : _GEN_257; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_259 = 9'h103 == io_addr ? mem_259 : _GEN_258; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_260 = 9'h104 == io_addr ? mem_260 : _GEN_259; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_261 = 9'h105 == io_addr ? mem_261 : _GEN_260; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_262 = 9'h106 == io_addr ? mem_262 : _GEN_261; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_263 = 9'h107 == io_addr ? mem_263 : _GEN_262; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_264 = 9'h108 == io_addr ? mem_264 : _GEN_263; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_265 = 9'h109 == io_addr ? mem_265 : _GEN_264; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_266 = 9'h10a == io_addr ? mem_266 : _GEN_265; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_267 = 9'h10b == io_addr ? mem_267 : _GEN_266; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_268 = 9'h10c == io_addr ? mem_268 : _GEN_267; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_269 = 9'h10d == io_addr ? mem_269 : _GEN_268; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_270 = 9'h10e == io_addr ? mem_270 : _GEN_269; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_271 = 9'h10f == io_addr ? mem_271 : _GEN_270; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_272 = 9'h110 == io_addr ? mem_272 : _GEN_271; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_273 = 9'h111 == io_addr ? mem_273 : _GEN_272; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_274 = 9'h112 == io_addr ? mem_274 : _GEN_273; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_275 = 9'h113 == io_addr ? mem_275 : _GEN_274; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_276 = 9'h114 == io_addr ? mem_276 : _GEN_275; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_277 = 9'h115 == io_addr ? mem_277 : _GEN_276; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_278 = 9'h116 == io_addr ? mem_278 : _GEN_277; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_279 = 9'h117 == io_addr ? mem_279 : _GEN_278; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_280 = 9'h118 == io_addr ? mem_280 : _GEN_279; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_281 = 9'h119 == io_addr ? mem_281 : _GEN_280; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_282 = 9'h11a == io_addr ? mem_282 : _GEN_281; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_283 = 9'h11b == io_addr ? mem_283 : _GEN_282; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_284 = 9'h11c == io_addr ? mem_284 : _GEN_283; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_285 = 9'h11d == io_addr ? mem_285 : _GEN_284; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_286 = 9'h11e == io_addr ? mem_286 : _GEN_285; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_287 = 9'h11f == io_addr ? mem_287 : _GEN_286; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_288 = 9'h120 == io_addr ? mem_288 : _GEN_287; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_289 = 9'h121 == io_addr ? mem_289 : _GEN_288; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_290 = 9'h122 == io_addr ? mem_290 : _GEN_289; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_291 = 9'h123 == io_addr ? mem_291 : _GEN_290; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_292 = 9'h124 == io_addr ? mem_292 : _GEN_291; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_293 = 9'h125 == io_addr ? mem_293 : _GEN_292; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_294 = 9'h126 == io_addr ? mem_294 : _GEN_293; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_295 = 9'h127 == io_addr ? mem_295 : _GEN_294; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_296 = 9'h128 == io_addr ? mem_296 : _GEN_295; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_297 = 9'h129 == io_addr ? mem_297 : _GEN_296; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_298 = 9'h12a == io_addr ? mem_298 : _GEN_297; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_299 = 9'h12b == io_addr ? mem_299 : _GEN_298; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_300 = 9'h12c == io_addr ? mem_300 : _GEN_299; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_301 = 9'h12d == io_addr ? mem_301 : _GEN_300; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_302 = 9'h12e == io_addr ? mem_302 : _GEN_301; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_303 = 9'h12f == io_addr ? mem_303 : _GEN_302; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_304 = 9'h130 == io_addr ? mem_304 : _GEN_303; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_305 = 9'h131 == io_addr ? mem_305 : _GEN_304; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_306 = 9'h132 == io_addr ? mem_306 : _GEN_305; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_307 = 9'h133 == io_addr ? mem_307 : _GEN_306; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_308 = 9'h134 == io_addr ? mem_308 : _GEN_307; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_309 = 9'h135 == io_addr ? mem_309 : _GEN_308; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_310 = 9'h136 == io_addr ? mem_310 : _GEN_309; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_311 = 9'h137 == io_addr ? mem_311 : _GEN_310; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_312 = 9'h138 == io_addr ? mem_312 : _GEN_311; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_313 = 9'h139 == io_addr ? mem_313 : _GEN_312; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_314 = 9'h13a == io_addr ? mem_314 : _GEN_313; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_315 = 9'h13b == io_addr ? mem_315 : _GEN_314; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_316 = 9'h13c == io_addr ? mem_316 : _GEN_315; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_317 = 9'h13d == io_addr ? mem_317 : _GEN_316; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_318 = 9'h13e == io_addr ? mem_318 : _GEN_317; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_319 = 9'h13f == io_addr ? mem_319 : _GEN_318; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_320 = 9'h140 == io_addr ? mem_320 : _GEN_319; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_321 = 9'h141 == io_addr ? mem_321 : _GEN_320; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_322 = 9'h142 == io_addr ? mem_322 : _GEN_321; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_323 = 9'h143 == io_addr ? mem_323 : _GEN_322; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_324 = 9'h144 == io_addr ? mem_324 : _GEN_323; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_325 = 9'h145 == io_addr ? mem_325 : _GEN_324; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_326 = 9'h146 == io_addr ? mem_326 : _GEN_325; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_327 = 9'h147 == io_addr ? mem_327 : _GEN_326; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_328 = 9'h148 == io_addr ? mem_328 : _GEN_327; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_329 = 9'h149 == io_addr ? mem_329 : _GEN_328; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_330 = 9'h14a == io_addr ? mem_330 : _GEN_329; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_331 = 9'h14b == io_addr ? mem_331 : _GEN_330; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_332 = 9'h14c == io_addr ? mem_332 : _GEN_331; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_333 = 9'h14d == io_addr ? mem_333 : _GEN_332; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_334 = 9'h14e == io_addr ? mem_334 : _GEN_333; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_335 = 9'h14f == io_addr ? mem_335 : _GEN_334; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_336 = 9'h150 == io_addr ? mem_336 : _GEN_335; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_337 = 9'h151 == io_addr ? mem_337 : _GEN_336; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_338 = 9'h152 == io_addr ? mem_338 : _GEN_337; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_339 = 9'h153 == io_addr ? mem_339 : _GEN_338; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_340 = 9'h154 == io_addr ? mem_340 : _GEN_339; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_341 = 9'h155 == io_addr ? mem_341 : _GEN_340; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_342 = 9'h156 == io_addr ? mem_342 : _GEN_341; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_343 = 9'h157 == io_addr ? mem_343 : _GEN_342; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_344 = 9'h158 == io_addr ? mem_344 : _GEN_343; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_345 = 9'h159 == io_addr ? mem_345 : _GEN_344; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_346 = 9'h15a == io_addr ? mem_346 : _GEN_345; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_347 = 9'h15b == io_addr ? mem_347 : _GEN_346; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_348 = 9'h15c == io_addr ? mem_348 : _GEN_347; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_349 = 9'h15d == io_addr ? mem_349 : _GEN_348; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_350 = 9'h15e == io_addr ? mem_350 : _GEN_349; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_351 = 9'h15f == io_addr ? mem_351 : _GEN_350; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_352 = 9'h160 == io_addr ? mem_352 : _GEN_351; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_353 = 9'h161 == io_addr ? mem_353 : _GEN_352; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_354 = 9'h162 == io_addr ? mem_354 : _GEN_353; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_355 = 9'h163 == io_addr ? mem_355 : _GEN_354; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_356 = 9'h164 == io_addr ? mem_356 : _GEN_355; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_357 = 9'h165 == io_addr ? mem_357 : _GEN_356; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_358 = 9'h166 == io_addr ? mem_358 : _GEN_357; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_359 = 9'h167 == io_addr ? mem_359 : _GEN_358; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_360 = 9'h168 == io_addr ? mem_360 : _GEN_359; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_361 = 9'h169 == io_addr ? mem_361 : _GEN_360; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_362 = 9'h16a == io_addr ? mem_362 : _GEN_361; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_363 = 9'h16b == io_addr ? mem_363 : _GEN_362; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_364 = 9'h16c == io_addr ? mem_364 : _GEN_363; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_365 = 9'h16d == io_addr ? mem_365 : _GEN_364; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_366 = 9'h16e == io_addr ? mem_366 : _GEN_365; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_367 = 9'h16f == io_addr ? mem_367 : _GEN_366; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_368 = 9'h170 == io_addr ? mem_368 : _GEN_367; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_369 = 9'h171 == io_addr ? mem_369 : _GEN_368; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_370 = 9'h172 == io_addr ? mem_370 : _GEN_369; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_371 = 9'h173 == io_addr ? mem_371 : _GEN_370; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_372 = 9'h174 == io_addr ? mem_372 : _GEN_371; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_373 = 9'h175 == io_addr ? mem_373 : _GEN_372; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_374 = 9'h176 == io_addr ? mem_374 : _GEN_373; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_375 = 9'h177 == io_addr ? mem_375 : _GEN_374; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_376 = 9'h178 == io_addr ? mem_376 : _GEN_375; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_377 = 9'h179 == io_addr ? mem_377 : _GEN_376; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_378 = 9'h17a == io_addr ? mem_378 : _GEN_377; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_379 = 9'h17b == io_addr ? mem_379 : _GEN_378; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_380 = 9'h17c == io_addr ? mem_380 : _GEN_379; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_381 = 9'h17d == io_addr ? mem_381 : _GEN_380; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_382 = 9'h17e == io_addr ? mem_382 : _GEN_381; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_383 = 9'h17f == io_addr ? mem_383 : _GEN_382; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_384 = 9'h180 == io_addr ? mem_384 : _GEN_383; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_385 = 9'h181 == io_addr ? mem_385 : _GEN_384; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_386 = 9'h182 == io_addr ? mem_386 : _GEN_385; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_387 = 9'h183 == io_addr ? mem_387 : _GEN_386; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_388 = 9'h184 == io_addr ? mem_388 : _GEN_387; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_389 = 9'h185 == io_addr ? mem_389 : _GEN_388; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_390 = 9'h186 == io_addr ? mem_390 : _GEN_389; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_391 = 9'h187 == io_addr ? mem_391 : _GEN_390; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_392 = 9'h188 == io_addr ? mem_392 : _GEN_391; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_393 = 9'h189 == io_addr ? mem_393 : _GEN_392; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_394 = 9'h18a == io_addr ? mem_394 : _GEN_393; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_395 = 9'h18b == io_addr ? mem_395 : _GEN_394; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_396 = 9'h18c == io_addr ? mem_396 : _GEN_395; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_397 = 9'h18d == io_addr ? mem_397 : _GEN_396; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_398 = 9'h18e == io_addr ? mem_398 : _GEN_397; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_399 = 9'h18f == io_addr ? mem_399 : _GEN_398; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_400 = 9'h190 == io_addr ? mem_400 : _GEN_399; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_401 = 9'h191 == io_addr ? mem_401 : _GEN_400; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_402 = 9'h192 == io_addr ? mem_402 : _GEN_401; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_403 = 9'h193 == io_addr ? mem_403 : _GEN_402; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_404 = 9'h194 == io_addr ? mem_404 : _GEN_403; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_405 = 9'h195 == io_addr ? mem_405 : _GEN_404; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_406 = 9'h196 == io_addr ? mem_406 : _GEN_405; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_407 = 9'h197 == io_addr ? mem_407 : _GEN_406; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_408 = 9'h198 == io_addr ? mem_408 : _GEN_407; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_409 = 9'h199 == io_addr ? mem_409 : _GEN_408; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_410 = 9'h19a == io_addr ? mem_410 : _GEN_409; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_411 = 9'h19b == io_addr ? mem_411 : _GEN_410; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_412 = 9'h19c == io_addr ? mem_412 : _GEN_411; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_413 = 9'h19d == io_addr ? mem_413 : _GEN_412; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_414 = 9'h19e == io_addr ? mem_414 : _GEN_413; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_415 = 9'h19f == io_addr ? mem_415 : _GEN_414; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_416 = 9'h1a0 == io_addr ? mem_416 : _GEN_415; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_417 = 9'h1a1 == io_addr ? mem_417 : _GEN_416; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_418 = 9'h1a2 == io_addr ? mem_418 : _GEN_417; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_419 = 9'h1a3 == io_addr ? mem_419 : _GEN_418; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_420 = 9'h1a4 == io_addr ? mem_420 : _GEN_419; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_421 = 9'h1a5 == io_addr ? mem_421 : _GEN_420; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_422 = 9'h1a6 == io_addr ? mem_422 : _GEN_421; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_423 = 9'h1a7 == io_addr ? mem_423 : _GEN_422; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_424 = 9'h1a8 == io_addr ? mem_424 : _GEN_423; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_425 = 9'h1a9 == io_addr ? mem_425 : _GEN_424; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_426 = 9'h1aa == io_addr ? mem_426 : _GEN_425; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_427 = 9'h1ab == io_addr ? mem_427 : _GEN_426; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_428 = 9'h1ac == io_addr ? mem_428 : _GEN_427; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_429 = 9'h1ad == io_addr ? mem_429 : _GEN_428; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_430 = 9'h1ae == io_addr ? mem_430 : _GEN_429; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_431 = 9'h1af == io_addr ? mem_431 : _GEN_430; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_432 = 9'h1b0 == io_addr ? mem_432 : _GEN_431; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_433 = 9'h1b1 == io_addr ? mem_433 : _GEN_432; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_434 = 9'h1b2 == io_addr ? mem_434 : _GEN_433; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_435 = 9'h1b3 == io_addr ? mem_435 : _GEN_434; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_436 = 9'h1b4 == io_addr ? mem_436 : _GEN_435; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_437 = 9'h1b5 == io_addr ? mem_437 : _GEN_436; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_438 = 9'h1b6 == io_addr ? mem_438 : _GEN_437; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_439 = 9'h1b7 == io_addr ? mem_439 : _GEN_438; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_440 = 9'h1b8 == io_addr ? mem_440 : _GEN_439; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_441 = 9'h1b9 == io_addr ? mem_441 : _GEN_440; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_442 = 9'h1ba == io_addr ? mem_442 : _GEN_441; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_443 = 9'h1bb == io_addr ? mem_443 : _GEN_442; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_444 = 9'h1bc == io_addr ? mem_444 : _GEN_443; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_445 = 9'h1bd == io_addr ? mem_445 : _GEN_444; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_446 = 9'h1be == io_addr ? mem_446 : _GEN_445; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_447 = 9'h1bf == io_addr ? mem_447 : _GEN_446; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_448 = 9'h1c0 == io_addr ? mem_448 : _GEN_447; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_449 = 9'h1c1 == io_addr ? mem_449 : _GEN_448; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_450 = 9'h1c2 == io_addr ? mem_450 : _GEN_449; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_451 = 9'h1c3 == io_addr ? mem_451 : _GEN_450; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_452 = 9'h1c4 == io_addr ? mem_452 : _GEN_451; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_453 = 9'h1c5 == io_addr ? mem_453 : _GEN_452; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_454 = 9'h1c6 == io_addr ? mem_454 : _GEN_453; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_455 = 9'h1c7 == io_addr ? mem_455 : _GEN_454; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_456 = 9'h1c8 == io_addr ? mem_456 : _GEN_455; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_457 = 9'h1c9 == io_addr ? mem_457 : _GEN_456; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_458 = 9'h1ca == io_addr ? mem_458 : _GEN_457; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_459 = 9'h1cb == io_addr ? mem_459 : _GEN_458; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_460 = 9'h1cc == io_addr ? mem_460 : _GEN_459; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_461 = 9'h1cd == io_addr ? mem_461 : _GEN_460; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_462 = 9'h1ce == io_addr ? mem_462 : _GEN_461; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_463 = 9'h1cf == io_addr ? mem_463 : _GEN_462; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_464 = 9'h1d0 == io_addr ? mem_464 : _GEN_463; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_465 = 9'h1d1 == io_addr ? mem_465 : _GEN_464; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_466 = 9'h1d2 == io_addr ? mem_466 : _GEN_465; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_467 = 9'h1d3 == io_addr ? mem_467 : _GEN_466; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_468 = 9'h1d4 == io_addr ? mem_468 : _GEN_467; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_469 = 9'h1d5 == io_addr ? mem_469 : _GEN_468; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_470 = 9'h1d6 == io_addr ? mem_470 : _GEN_469; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_471 = 9'h1d7 == io_addr ? mem_471 : _GEN_470; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_472 = 9'h1d8 == io_addr ? mem_472 : _GEN_471; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_473 = 9'h1d9 == io_addr ? mem_473 : _GEN_472; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_474 = 9'h1da == io_addr ? mem_474 : _GEN_473; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_475 = 9'h1db == io_addr ? mem_475 : _GEN_474; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_476 = 9'h1dc == io_addr ? mem_476 : _GEN_475; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_477 = 9'h1dd == io_addr ? mem_477 : _GEN_476; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_478 = 9'h1de == io_addr ? mem_478 : _GEN_477; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_479 = 9'h1df == io_addr ? mem_479 : _GEN_478; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_480 = 9'h1e0 == io_addr ? mem_480 : _GEN_479; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_481 = 9'h1e1 == io_addr ? mem_481 : _GEN_480; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_482 = 9'h1e2 == io_addr ? mem_482 : _GEN_481; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_483 = 9'h1e3 == io_addr ? mem_483 : _GEN_482; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_484 = 9'h1e4 == io_addr ? mem_484 : _GEN_483; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_485 = 9'h1e5 == io_addr ? mem_485 : _GEN_484; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_486 = 9'h1e6 == io_addr ? mem_486 : _GEN_485; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_487 = 9'h1e7 == io_addr ? mem_487 : _GEN_486; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_488 = 9'h1e8 == io_addr ? mem_488 : _GEN_487; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_489 = 9'h1e9 == io_addr ? mem_489 : _GEN_488; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_490 = 9'h1ea == io_addr ? mem_490 : _GEN_489; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_491 = 9'h1eb == io_addr ? mem_491 : _GEN_490; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_492 = 9'h1ec == io_addr ? mem_492 : _GEN_491; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_493 = 9'h1ed == io_addr ? mem_493 : _GEN_492; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_494 = 9'h1ee == io_addr ? mem_494 : _GEN_493; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_495 = 9'h1ef == io_addr ? mem_495 : _GEN_494; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_496 = 9'h1f0 == io_addr ? mem_496 : _GEN_495; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_497 = 9'h1f1 == io_addr ? mem_497 : _GEN_496; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_498 = 9'h1f2 == io_addr ? mem_498 : _GEN_497; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_499 = 9'h1f3 == io_addr ? mem_499 : _GEN_498; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_500 = 9'h1f4 == io_addr ? mem_500 : _GEN_499; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_501 = 9'h1f5 == io_addr ? mem_501 : _GEN_500; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_502 = 9'h1f6 == io_addr ? mem_502 : _GEN_501; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_503 = 9'h1f7 == io_addr ? mem_503 : _GEN_502; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_504 = 9'h1f8 == io_addr ? mem_504 : _GEN_503; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_505 = 9'h1f9 == io_addr ? mem_505 : _GEN_504; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_506 = 9'h1fa == io_addr ? mem_506 : _GEN_505; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [255:0] _GEN_507 = 9'h1fb == io_addr ? mem_507 : _GEN_506; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  assign io_dout = io_dout_REG; // @[RAMWrapper.scala 288:11]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_0 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_0 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_1 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_1 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_2 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_2 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_3 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_3 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_4 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_4 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_5 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_5 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_6 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_6 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_7 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_7 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_8 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_8 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_9 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_9 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_10 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_10 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_11 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_11 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_12 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_12 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_13 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_13 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_14 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_14 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_15 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_15 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_16 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_16 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_17 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_17 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_18 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_18 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_19 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_19 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_20 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_20 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_21 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_21 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_22 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_22 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_23 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_23 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_24 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_24 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_25 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_25 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_26 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_26 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_27 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_27 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_28 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_28 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_29 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_29 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_30 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_30 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_31 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_31 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_32 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h20 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_32 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_33 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h21 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_33 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_34 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h22 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_34 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_35 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h23 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_35 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_36 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h24 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_36 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_37 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h25 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_37 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_38 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h26 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_38 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_39 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h27 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_39 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_40 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h28 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_40 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_41 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h29 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_41 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_42 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_42 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_43 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_43 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_44 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_44 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_45 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_45 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_46 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_46 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_47 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_47 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_48 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h30 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_48 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_49 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h31 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_49 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_50 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h32 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_50 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_51 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h33 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_51 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_52 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h34 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_52 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_53 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h35 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_53 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_54 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h36 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_54 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_55 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h37 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_55 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_56 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h38 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_56 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_57 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h39 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_57 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_58 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_58 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_59 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_59 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_60 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_60 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_61 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_61 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_62 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_62 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_63 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_63 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_64 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h40 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_64 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_65 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h41 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_65 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_66 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h42 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_66 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_67 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h43 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_67 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_68 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h44 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_68 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_69 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h45 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_69 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_70 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h46 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_70 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_71 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h47 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_71 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_72 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h48 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_72 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_73 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h49 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_73 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_74 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_74 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_75 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_75 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_76 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_76 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_77 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_77 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_78 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_78 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_79 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_79 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_80 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h50 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_80 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_81 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h51 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_81 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_82 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h52 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_82 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_83 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h53 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_83 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_84 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h54 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_84 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_85 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h55 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_85 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_86 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h56 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_86 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_87 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h57 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_87 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_88 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h58 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_88 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_89 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h59 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_89 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_90 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_90 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_91 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_91 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_92 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_92 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_93 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_93 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_94 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_94 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_95 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_95 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_96 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h60 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_96 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_97 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h61 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_97 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_98 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h62 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_98 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_99 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h63 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_99 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_100 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h64 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_100 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_101 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h65 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_101 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_102 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h66 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_102 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_103 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h67 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_103 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_104 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h68 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_104 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_105 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h69 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_105 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_106 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_106 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_107 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_107 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_108 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_108 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_109 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_109 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_110 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_110 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_111 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_111 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_112 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h70 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_112 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_113 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h71 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_113 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_114 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h72 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_114 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_115 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h73 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_115 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_116 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h74 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_116 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_117 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h75 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_117 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_118 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h76 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_118 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_119 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h77 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_119 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_120 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h78 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_120 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_121 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h79 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_121 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_122 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_122 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_123 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_123 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_124 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_124 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_125 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_125 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_126 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_126 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_127 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_127 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_128 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h80 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_128 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_129 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h81 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_129 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_130 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h82 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_130 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_131 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h83 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_131 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_132 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h84 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_132 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_133 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h85 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_133 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_134 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h86 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_134 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_135 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h87 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_135 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_136 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h88 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_136 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_137 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h89 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_137 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_138 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_138 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_139 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_139 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_140 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_140 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_141 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_141 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_142 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_142 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_143 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_143 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_144 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h90 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_144 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_145 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h91 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_145 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_146 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h92 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_146 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_147 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h93 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_147 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_148 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h94 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_148 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_149 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h95 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_149 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_150 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h96 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_150 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_151 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h97 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_151 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_152 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h98 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_152 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_153 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h99 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_153 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_154 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_154 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_155 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_155 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_156 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_156 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_157 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_157 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_158 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_158 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_159 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_159 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_160 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_160 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_161 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_161 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_162 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_162 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_163 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_163 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_164 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_164 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_165 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_165 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_166 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_166 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_167 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_167 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_168 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_168 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_169 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_169 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_170 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'haa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_170 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_171 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hab == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_171 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_172 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hac == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_172 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_173 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'had == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_173 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_174 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hae == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_174 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_175 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'haf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_175 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_176 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_176 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_177 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_177 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_178 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_178 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_179 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_179 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_180 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_180 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_181 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_181 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_182 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_182 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_183 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_183 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_184 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_184 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_185 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_185 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_186 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hba == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_186 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_187 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_187 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_188 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_188 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_189 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_189 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_190 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_190 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_191 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_191 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_192 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_192 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_193 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_193 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_194 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_194 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_195 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_195 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_196 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_196 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_197 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_197 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_198 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_198 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_199 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_199 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_200 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_200 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_201 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_201 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_202 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hca == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_202 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_203 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_203 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_204 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_204 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_205 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_205 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_206 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hce == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_206 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_207 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_207 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_208 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_208 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_209 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_209 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_210 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_210 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_211 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_211 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_212 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_212 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_213 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_213 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_214 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_214 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_215 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_215 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_216 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_216 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_217 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_217 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_218 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hda == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_218 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_219 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_219 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_220 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_220 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_221 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_221 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_222 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hde == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_222 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_223 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_223 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_224 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_224 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_225 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_225 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_226 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_226 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_227 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_227 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_228 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_228 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_229 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_229 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_230 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_230 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_231 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_231 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_232 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_232 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_233 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_233 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_234 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hea == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_234 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_235 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'heb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_235 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_236 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hec == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_236 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_237 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hed == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_237 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_238 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hee == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_238 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_239 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hef == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_239 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_240 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_240 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_241 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_241 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_242 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_242 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_243 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_243 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_244 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_244 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_245 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_245 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_246 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_246 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_247 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_247 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_248 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_248 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_249 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_249 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_250 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_250 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_251 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_251 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_252 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_252 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_253 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_253 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_254 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_254 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_255 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hff == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_255 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_256 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h100 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_256 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_257 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h101 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_257 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_258 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h102 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_258 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_259 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h103 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_259 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_260 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h104 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_260 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_261 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h105 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_261 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_262 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h106 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_262 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_263 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h107 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_263 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_264 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h108 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_264 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_265 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h109 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_265 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_266 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_266 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_267 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_267 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_268 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_268 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_269 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_269 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_270 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_270 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_271 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_271 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_272 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h110 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_272 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_273 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h111 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_273 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_274 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h112 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_274 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_275 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h113 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_275 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_276 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h114 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_276 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_277 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h115 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_277 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_278 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h116 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_278 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_279 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h117 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_279 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_280 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h118 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_280 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_281 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h119 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_281 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_282 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_282 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_283 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_283 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_284 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_284 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_285 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_285 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_286 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_286 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_287 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_287 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_288 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h120 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_288 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_289 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h121 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_289 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_290 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h122 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_290 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_291 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h123 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_291 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_292 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h124 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_292 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_293 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h125 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_293 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_294 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h126 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_294 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_295 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h127 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_295 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_296 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h128 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_296 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_297 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h129 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_297 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_298 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_298 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_299 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_299 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_300 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_300 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_301 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_301 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_302 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_302 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_303 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_303 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_304 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h130 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_304 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_305 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h131 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_305 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_306 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h132 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_306 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_307 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h133 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_307 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_308 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h134 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_308 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_309 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h135 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_309 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_310 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h136 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_310 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_311 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h137 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_311 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_312 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h138 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_312 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_313 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h139 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_313 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_314 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_314 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_315 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_315 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_316 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_316 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_317 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_317 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_318 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_318 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_319 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_319 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_320 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h140 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_320 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_321 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h141 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_321 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_322 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h142 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_322 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_323 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h143 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_323 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_324 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h144 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_324 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_325 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h145 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_325 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_326 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h146 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_326 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_327 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h147 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_327 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_328 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h148 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_328 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_329 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h149 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_329 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_330 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_330 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_331 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_331 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_332 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_332 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_333 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_333 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_334 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_334 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_335 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_335 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_336 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h150 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_336 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_337 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h151 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_337 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_338 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h152 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_338 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_339 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h153 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_339 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_340 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h154 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_340 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_341 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h155 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_341 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_342 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h156 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_342 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_343 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h157 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_343 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_344 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h158 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_344 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_345 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h159 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_345 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_346 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_346 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_347 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_347 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_348 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_348 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_349 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_349 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_350 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_350 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_351 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_351 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_352 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h160 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_352 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_353 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h161 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_353 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_354 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h162 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_354 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_355 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h163 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_355 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_356 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h164 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_356 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_357 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h165 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_357 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_358 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h166 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_358 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_359 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h167 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_359 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_360 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h168 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_360 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_361 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h169 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_361 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_362 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_362 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_363 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_363 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_364 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_364 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_365 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_365 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_366 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_366 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_367 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_367 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_368 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h170 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_368 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_369 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h171 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_369 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_370 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h172 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_370 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_371 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h173 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_371 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_372 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h174 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_372 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_373 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h175 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_373 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_374 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h176 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_374 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_375 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h177 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_375 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_376 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h178 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_376 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_377 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h179 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_377 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_378 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_378 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_379 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_379 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_380 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_380 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_381 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_381 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_382 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_382 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_383 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_383 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_384 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h180 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_384 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_385 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h181 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_385 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_386 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h182 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_386 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_387 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h183 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_387 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_388 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h184 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_388 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_389 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h185 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_389 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_390 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h186 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_390 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_391 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h187 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_391 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_392 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h188 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_392 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_393 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h189 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_393 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_394 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_394 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_395 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_395 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_396 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_396 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_397 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_397 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_398 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_398 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_399 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_399 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_400 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h190 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_400 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_401 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h191 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_401 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_402 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h192 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_402 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_403 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h193 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_403 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_404 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h194 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_404 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_405 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h195 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_405 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_406 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h196 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_406 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_407 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h197 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_407 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_408 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h198 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_408 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_409 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h199 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_409 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_410 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_410 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_411 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_411 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_412 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_412 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_413 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_413 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_414 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_414 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_415 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_415 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_416 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_416 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_417 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_417 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_418 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_418 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_419 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_419 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_420 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_420 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_421 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_421 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_422 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_422 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_423 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_423 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_424 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_424 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_425 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_425 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_426 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1aa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_426 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_427 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ab == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_427 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_428 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ac == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_428 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_429 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ad == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_429 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_430 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ae == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_430 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_431 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1af == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_431 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_432 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_432 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_433 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_433 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_434 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_434 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_435 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_435 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_436 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_436 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_437 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_437 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_438 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_438 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_439 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_439 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_440 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_440 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_441 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_441 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_442 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ba == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_442 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_443 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_443 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_444 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_444 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_445 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_445 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_446 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1be == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_446 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_447 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_447 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_448 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_448 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_449 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_449 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_450 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_450 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_451 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_451 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_452 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_452 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_453 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_453 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_454 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_454 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_455 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_455 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_456 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_456 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_457 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_457 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_458 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ca == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_458 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_459 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_459 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_460 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_460 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_461 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_461 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_462 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ce == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_462 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_463 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_463 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_464 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_464 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_465 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_465 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_466 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_466 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_467 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_467 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_468 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_468 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_469 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_469 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_470 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_470 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_471 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_471 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_472 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_472 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_473 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_473 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_474 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1da == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_474 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_475 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1db == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_475 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_476 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1dc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_476 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_477 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1dd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_477 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_478 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1de == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_478 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_479 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1df == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_479 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_480 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_480 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_481 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_481 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_482 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_482 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_483 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_483 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_484 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_484 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_485 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_485 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_486 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_486 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_487 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_487 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_488 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_488 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_489 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_489 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_490 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ea == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_490 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_491 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1eb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_491 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_492 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ec == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_492 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_493 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ed == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_493 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_494 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ee == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_494 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_495 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ef == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_495 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_496 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_496 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_497 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_497 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_498 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_498 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_499 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_499 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_500 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_500 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_501 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_501 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_502 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_502 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_503 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_503 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_504 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_504 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_505 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_505 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_506 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_506 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_507 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_507 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_508 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_508 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_509 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_509 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_510 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_510 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_511 <= 256'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ff == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_511 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (9'h1ff == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_511; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fe == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_510; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fd == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_509; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fc == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_508; // @[RAMWrapper.scala 288:21]
    end else begin
      io_dout_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  mem_0 = _RAND_0[255:0];
  _RAND_1 = {8{`RANDOM}};
  mem_1 = _RAND_1[255:0];
  _RAND_2 = {8{`RANDOM}};
  mem_2 = _RAND_2[255:0];
  _RAND_3 = {8{`RANDOM}};
  mem_3 = _RAND_3[255:0];
  _RAND_4 = {8{`RANDOM}};
  mem_4 = _RAND_4[255:0];
  _RAND_5 = {8{`RANDOM}};
  mem_5 = _RAND_5[255:0];
  _RAND_6 = {8{`RANDOM}};
  mem_6 = _RAND_6[255:0];
  _RAND_7 = {8{`RANDOM}};
  mem_7 = _RAND_7[255:0];
  _RAND_8 = {8{`RANDOM}};
  mem_8 = _RAND_8[255:0];
  _RAND_9 = {8{`RANDOM}};
  mem_9 = _RAND_9[255:0];
  _RAND_10 = {8{`RANDOM}};
  mem_10 = _RAND_10[255:0];
  _RAND_11 = {8{`RANDOM}};
  mem_11 = _RAND_11[255:0];
  _RAND_12 = {8{`RANDOM}};
  mem_12 = _RAND_12[255:0];
  _RAND_13 = {8{`RANDOM}};
  mem_13 = _RAND_13[255:0];
  _RAND_14 = {8{`RANDOM}};
  mem_14 = _RAND_14[255:0];
  _RAND_15 = {8{`RANDOM}};
  mem_15 = _RAND_15[255:0];
  _RAND_16 = {8{`RANDOM}};
  mem_16 = _RAND_16[255:0];
  _RAND_17 = {8{`RANDOM}};
  mem_17 = _RAND_17[255:0];
  _RAND_18 = {8{`RANDOM}};
  mem_18 = _RAND_18[255:0];
  _RAND_19 = {8{`RANDOM}};
  mem_19 = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  mem_20 = _RAND_20[255:0];
  _RAND_21 = {8{`RANDOM}};
  mem_21 = _RAND_21[255:0];
  _RAND_22 = {8{`RANDOM}};
  mem_22 = _RAND_22[255:0];
  _RAND_23 = {8{`RANDOM}};
  mem_23 = _RAND_23[255:0];
  _RAND_24 = {8{`RANDOM}};
  mem_24 = _RAND_24[255:0];
  _RAND_25 = {8{`RANDOM}};
  mem_25 = _RAND_25[255:0];
  _RAND_26 = {8{`RANDOM}};
  mem_26 = _RAND_26[255:0];
  _RAND_27 = {8{`RANDOM}};
  mem_27 = _RAND_27[255:0];
  _RAND_28 = {8{`RANDOM}};
  mem_28 = _RAND_28[255:0];
  _RAND_29 = {8{`RANDOM}};
  mem_29 = _RAND_29[255:0];
  _RAND_30 = {8{`RANDOM}};
  mem_30 = _RAND_30[255:0];
  _RAND_31 = {8{`RANDOM}};
  mem_31 = _RAND_31[255:0];
  _RAND_32 = {8{`RANDOM}};
  mem_32 = _RAND_32[255:0];
  _RAND_33 = {8{`RANDOM}};
  mem_33 = _RAND_33[255:0];
  _RAND_34 = {8{`RANDOM}};
  mem_34 = _RAND_34[255:0];
  _RAND_35 = {8{`RANDOM}};
  mem_35 = _RAND_35[255:0];
  _RAND_36 = {8{`RANDOM}};
  mem_36 = _RAND_36[255:0];
  _RAND_37 = {8{`RANDOM}};
  mem_37 = _RAND_37[255:0];
  _RAND_38 = {8{`RANDOM}};
  mem_38 = _RAND_38[255:0];
  _RAND_39 = {8{`RANDOM}};
  mem_39 = _RAND_39[255:0];
  _RAND_40 = {8{`RANDOM}};
  mem_40 = _RAND_40[255:0];
  _RAND_41 = {8{`RANDOM}};
  mem_41 = _RAND_41[255:0];
  _RAND_42 = {8{`RANDOM}};
  mem_42 = _RAND_42[255:0];
  _RAND_43 = {8{`RANDOM}};
  mem_43 = _RAND_43[255:0];
  _RAND_44 = {8{`RANDOM}};
  mem_44 = _RAND_44[255:0];
  _RAND_45 = {8{`RANDOM}};
  mem_45 = _RAND_45[255:0];
  _RAND_46 = {8{`RANDOM}};
  mem_46 = _RAND_46[255:0];
  _RAND_47 = {8{`RANDOM}};
  mem_47 = _RAND_47[255:0];
  _RAND_48 = {8{`RANDOM}};
  mem_48 = _RAND_48[255:0];
  _RAND_49 = {8{`RANDOM}};
  mem_49 = _RAND_49[255:0];
  _RAND_50 = {8{`RANDOM}};
  mem_50 = _RAND_50[255:0];
  _RAND_51 = {8{`RANDOM}};
  mem_51 = _RAND_51[255:0];
  _RAND_52 = {8{`RANDOM}};
  mem_52 = _RAND_52[255:0];
  _RAND_53 = {8{`RANDOM}};
  mem_53 = _RAND_53[255:0];
  _RAND_54 = {8{`RANDOM}};
  mem_54 = _RAND_54[255:0];
  _RAND_55 = {8{`RANDOM}};
  mem_55 = _RAND_55[255:0];
  _RAND_56 = {8{`RANDOM}};
  mem_56 = _RAND_56[255:0];
  _RAND_57 = {8{`RANDOM}};
  mem_57 = _RAND_57[255:0];
  _RAND_58 = {8{`RANDOM}};
  mem_58 = _RAND_58[255:0];
  _RAND_59 = {8{`RANDOM}};
  mem_59 = _RAND_59[255:0];
  _RAND_60 = {8{`RANDOM}};
  mem_60 = _RAND_60[255:0];
  _RAND_61 = {8{`RANDOM}};
  mem_61 = _RAND_61[255:0];
  _RAND_62 = {8{`RANDOM}};
  mem_62 = _RAND_62[255:0];
  _RAND_63 = {8{`RANDOM}};
  mem_63 = _RAND_63[255:0];
  _RAND_64 = {8{`RANDOM}};
  mem_64 = _RAND_64[255:0];
  _RAND_65 = {8{`RANDOM}};
  mem_65 = _RAND_65[255:0];
  _RAND_66 = {8{`RANDOM}};
  mem_66 = _RAND_66[255:0];
  _RAND_67 = {8{`RANDOM}};
  mem_67 = _RAND_67[255:0];
  _RAND_68 = {8{`RANDOM}};
  mem_68 = _RAND_68[255:0];
  _RAND_69 = {8{`RANDOM}};
  mem_69 = _RAND_69[255:0];
  _RAND_70 = {8{`RANDOM}};
  mem_70 = _RAND_70[255:0];
  _RAND_71 = {8{`RANDOM}};
  mem_71 = _RAND_71[255:0];
  _RAND_72 = {8{`RANDOM}};
  mem_72 = _RAND_72[255:0];
  _RAND_73 = {8{`RANDOM}};
  mem_73 = _RAND_73[255:0];
  _RAND_74 = {8{`RANDOM}};
  mem_74 = _RAND_74[255:0];
  _RAND_75 = {8{`RANDOM}};
  mem_75 = _RAND_75[255:0];
  _RAND_76 = {8{`RANDOM}};
  mem_76 = _RAND_76[255:0];
  _RAND_77 = {8{`RANDOM}};
  mem_77 = _RAND_77[255:0];
  _RAND_78 = {8{`RANDOM}};
  mem_78 = _RAND_78[255:0];
  _RAND_79 = {8{`RANDOM}};
  mem_79 = _RAND_79[255:0];
  _RAND_80 = {8{`RANDOM}};
  mem_80 = _RAND_80[255:0];
  _RAND_81 = {8{`RANDOM}};
  mem_81 = _RAND_81[255:0];
  _RAND_82 = {8{`RANDOM}};
  mem_82 = _RAND_82[255:0];
  _RAND_83 = {8{`RANDOM}};
  mem_83 = _RAND_83[255:0];
  _RAND_84 = {8{`RANDOM}};
  mem_84 = _RAND_84[255:0];
  _RAND_85 = {8{`RANDOM}};
  mem_85 = _RAND_85[255:0];
  _RAND_86 = {8{`RANDOM}};
  mem_86 = _RAND_86[255:0];
  _RAND_87 = {8{`RANDOM}};
  mem_87 = _RAND_87[255:0];
  _RAND_88 = {8{`RANDOM}};
  mem_88 = _RAND_88[255:0];
  _RAND_89 = {8{`RANDOM}};
  mem_89 = _RAND_89[255:0];
  _RAND_90 = {8{`RANDOM}};
  mem_90 = _RAND_90[255:0];
  _RAND_91 = {8{`RANDOM}};
  mem_91 = _RAND_91[255:0];
  _RAND_92 = {8{`RANDOM}};
  mem_92 = _RAND_92[255:0];
  _RAND_93 = {8{`RANDOM}};
  mem_93 = _RAND_93[255:0];
  _RAND_94 = {8{`RANDOM}};
  mem_94 = _RAND_94[255:0];
  _RAND_95 = {8{`RANDOM}};
  mem_95 = _RAND_95[255:0];
  _RAND_96 = {8{`RANDOM}};
  mem_96 = _RAND_96[255:0];
  _RAND_97 = {8{`RANDOM}};
  mem_97 = _RAND_97[255:0];
  _RAND_98 = {8{`RANDOM}};
  mem_98 = _RAND_98[255:0];
  _RAND_99 = {8{`RANDOM}};
  mem_99 = _RAND_99[255:0];
  _RAND_100 = {8{`RANDOM}};
  mem_100 = _RAND_100[255:0];
  _RAND_101 = {8{`RANDOM}};
  mem_101 = _RAND_101[255:0];
  _RAND_102 = {8{`RANDOM}};
  mem_102 = _RAND_102[255:0];
  _RAND_103 = {8{`RANDOM}};
  mem_103 = _RAND_103[255:0];
  _RAND_104 = {8{`RANDOM}};
  mem_104 = _RAND_104[255:0];
  _RAND_105 = {8{`RANDOM}};
  mem_105 = _RAND_105[255:0];
  _RAND_106 = {8{`RANDOM}};
  mem_106 = _RAND_106[255:0];
  _RAND_107 = {8{`RANDOM}};
  mem_107 = _RAND_107[255:0];
  _RAND_108 = {8{`RANDOM}};
  mem_108 = _RAND_108[255:0];
  _RAND_109 = {8{`RANDOM}};
  mem_109 = _RAND_109[255:0];
  _RAND_110 = {8{`RANDOM}};
  mem_110 = _RAND_110[255:0];
  _RAND_111 = {8{`RANDOM}};
  mem_111 = _RAND_111[255:0];
  _RAND_112 = {8{`RANDOM}};
  mem_112 = _RAND_112[255:0];
  _RAND_113 = {8{`RANDOM}};
  mem_113 = _RAND_113[255:0];
  _RAND_114 = {8{`RANDOM}};
  mem_114 = _RAND_114[255:0];
  _RAND_115 = {8{`RANDOM}};
  mem_115 = _RAND_115[255:0];
  _RAND_116 = {8{`RANDOM}};
  mem_116 = _RAND_116[255:0];
  _RAND_117 = {8{`RANDOM}};
  mem_117 = _RAND_117[255:0];
  _RAND_118 = {8{`RANDOM}};
  mem_118 = _RAND_118[255:0];
  _RAND_119 = {8{`RANDOM}};
  mem_119 = _RAND_119[255:0];
  _RAND_120 = {8{`RANDOM}};
  mem_120 = _RAND_120[255:0];
  _RAND_121 = {8{`RANDOM}};
  mem_121 = _RAND_121[255:0];
  _RAND_122 = {8{`RANDOM}};
  mem_122 = _RAND_122[255:0];
  _RAND_123 = {8{`RANDOM}};
  mem_123 = _RAND_123[255:0];
  _RAND_124 = {8{`RANDOM}};
  mem_124 = _RAND_124[255:0];
  _RAND_125 = {8{`RANDOM}};
  mem_125 = _RAND_125[255:0];
  _RAND_126 = {8{`RANDOM}};
  mem_126 = _RAND_126[255:0];
  _RAND_127 = {8{`RANDOM}};
  mem_127 = _RAND_127[255:0];
  _RAND_128 = {8{`RANDOM}};
  mem_128 = _RAND_128[255:0];
  _RAND_129 = {8{`RANDOM}};
  mem_129 = _RAND_129[255:0];
  _RAND_130 = {8{`RANDOM}};
  mem_130 = _RAND_130[255:0];
  _RAND_131 = {8{`RANDOM}};
  mem_131 = _RAND_131[255:0];
  _RAND_132 = {8{`RANDOM}};
  mem_132 = _RAND_132[255:0];
  _RAND_133 = {8{`RANDOM}};
  mem_133 = _RAND_133[255:0];
  _RAND_134 = {8{`RANDOM}};
  mem_134 = _RAND_134[255:0];
  _RAND_135 = {8{`RANDOM}};
  mem_135 = _RAND_135[255:0];
  _RAND_136 = {8{`RANDOM}};
  mem_136 = _RAND_136[255:0];
  _RAND_137 = {8{`RANDOM}};
  mem_137 = _RAND_137[255:0];
  _RAND_138 = {8{`RANDOM}};
  mem_138 = _RAND_138[255:0];
  _RAND_139 = {8{`RANDOM}};
  mem_139 = _RAND_139[255:0];
  _RAND_140 = {8{`RANDOM}};
  mem_140 = _RAND_140[255:0];
  _RAND_141 = {8{`RANDOM}};
  mem_141 = _RAND_141[255:0];
  _RAND_142 = {8{`RANDOM}};
  mem_142 = _RAND_142[255:0];
  _RAND_143 = {8{`RANDOM}};
  mem_143 = _RAND_143[255:0];
  _RAND_144 = {8{`RANDOM}};
  mem_144 = _RAND_144[255:0];
  _RAND_145 = {8{`RANDOM}};
  mem_145 = _RAND_145[255:0];
  _RAND_146 = {8{`RANDOM}};
  mem_146 = _RAND_146[255:0];
  _RAND_147 = {8{`RANDOM}};
  mem_147 = _RAND_147[255:0];
  _RAND_148 = {8{`RANDOM}};
  mem_148 = _RAND_148[255:0];
  _RAND_149 = {8{`RANDOM}};
  mem_149 = _RAND_149[255:0];
  _RAND_150 = {8{`RANDOM}};
  mem_150 = _RAND_150[255:0];
  _RAND_151 = {8{`RANDOM}};
  mem_151 = _RAND_151[255:0];
  _RAND_152 = {8{`RANDOM}};
  mem_152 = _RAND_152[255:0];
  _RAND_153 = {8{`RANDOM}};
  mem_153 = _RAND_153[255:0];
  _RAND_154 = {8{`RANDOM}};
  mem_154 = _RAND_154[255:0];
  _RAND_155 = {8{`RANDOM}};
  mem_155 = _RAND_155[255:0];
  _RAND_156 = {8{`RANDOM}};
  mem_156 = _RAND_156[255:0];
  _RAND_157 = {8{`RANDOM}};
  mem_157 = _RAND_157[255:0];
  _RAND_158 = {8{`RANDOM}};
  mem_158 = _RAND_158[255:0];
  _RAND_159 = {8{`RANDOM}};
  mem_159 = _RAND_159[255:0];
  _RAND_160 = {8{`RANDOM}};
  mem_160 = _RAND_160[255:0];
  _RAND_161 = {8{`RANDOM}};
  mem_161 = _RAND_161[255:0];
  _RAND_162 = {8{`RANDOM}};
  mem_162 = _RAND_162[255:0];
  _RAND_163 = {8{`RANDOM}};
  mem_163 = _RAND_163[255:0];
  _RAND_164 = {8{`RANDOM}};
  mem_164 = _RAND_164[255:0];
  _RAND_165 = {8{`RANDOM}};
  mem_165 = _RAND_165[255:0];
  _RAND_166 = {8{`RANDOM}};
  mem_166 = _RAND_166[255:0];
  _RAND_167 = {8{`RANDOM}};
  mem_167 = _RAND_167[255:0];
  _RAND_168 = {8{`RANDOM}};
  mem_168 = _RAND_168[255:0];
  _RAND_169 = {8{`RANDOM}};
  mem_169 = _RAND_169[255:0];
  _RAND_170 = {8{`RANDOM}};
  mem_170 = _RAND_170[255:0];
  _RAND_171 = {8{`RANDOM}};
  mem_171 = _RAND_171[255:0];
  _RAND_172 = {8{`RANDOM}};
  mem_172 = _RAND_172[255:0];
  _RAND_173 = {8{`RANDOM}};
  mem_173 = _RAND_173[255:0];
  _RAND_174 = {8{`RANDOM}};
  mem_174 = _RAND_174[255:0];
  _RAND_175 = {8{`RANDOM}};
  mem_175 = _RAND_175[255:0];
  _RAND_176 = {8{`RANDOM}};
  mem_176 = _RAND_176[255:0];
  _RAND_177 = {8{`RANDOM}};
  mem_177 = _RAND_177[255:0];
  _RAND_178 = {8{`RANDOM}};
  mem_178 = _RAND_178[255:0];
  _RAND_179 = {8{`RANDOM}};
  mem_179 = _RAND_179[255:0];
  _RAND_180 = {8{`RANDOM}};
  mem_180 = _RAND_180[255:0];
  _RAND_181 = {8{`RANDOM}};
  mem_181 = _RAND_181[255:0];
  _RAND_182 = {8{`RANDOM}};
  mem_182 = _RAND_182[255:0];
  _RAND_183 = {8{`RANDOM}};
  mem_183 = _RAND_183[255:0];
  _RAND_184 = {8{`RANDOM}};
  mem_184 = _RAND_184[255:0];
  _RAND_185 = {8{`RANDOM}};
  mem_185 = _RAND_185[255:0];
  _RAND_186 = {8{`RANDOM}};
  mem_186 = _RAND_186[255:0];
  _RAND_187 = {8{`RANDOM}};
  mem_187 = _RAND_187[255:0];
  _RAND_188 = {8{`RANDOM}};
  mem_188 = _RAND_188[255:0];
  _RAND_189 = {8{`RANDOM}};
  mem_189 = _RAND_189[255:0];
  _RAND_190 = {8{`RANDOM}};
  mem_190 = _RAND_190[255:0];
  _RAND_191 = {8{`RANDOM}};
  mem_191 = _RAND_191[255:0];
  _RAND_192 = {8{`RANDOM}};
  mem_192 = _RAND_192[255:0];
  _RAND_193 = {8{`RANDOM}};
  mem_193 = _RAND_193[255:0];
  _RAND_194 = {8{`RANDOM}};
  mem_194 = _RAND_194[255:0];
  _RAND_195 = {8{`RANDOM}};
  mem_195 = _RAND_195[255:0];
  _RAND_196 = {8{`RANDOM}};
  mem_196 = _RAND_196[255:0];
  _RAND_197 = {8{`RANDOM}};
  mem_197 = _RAND_197[255:0];
  _RAND_198 = {8{`RANDOM}};
  mem_198 = _RAND_198[255:0];
  _RAND_199 = {8{`RANDOM}};
  mem_199 = _RAND_199[255:0];
  _RAND_200 = {8{`RANDOM}};
  mem_200 = _RAND_200[255:0];
  _RAND_201 = {8{`RANDOM}};
  mem_201 = _RAND_201[255:0];
  _RAND_202 = {8{`RANDOM}};
  mem_202 = _RAND_202[255:0];
  _RAND_203 = {8{`RANDOM}};
  mem_203 = _RAND_203[255:0];
  _RAND_204 = {8{`RANDOM}};
  mem_204 = _RAND_204[255:0];
  _RAND_205 = {8{`RANDOM}};
  mem_205 = _RAND_205[255:0];
  _RAND_206 = {8{`RANDOM}};
  mem_206 = _RAND_206[255:0];
  _RAND_207 = {8{`RANDOM}};
  mem_207 = _RAND_207[255:0];
  _RAND_208 = {8{`RANDOM}};
  mem_208 = _RAND_208[255:0];
  _RAND_209 = {8{`RANDOM}};
  mem_209 = _RAND_209[255:0];
  _RAND_210 = {8{`RANDOM}};
  mem_210 = _RAND_210[255:0];
  _RAND_211 = {8{`RANDOM}};
  mem_211 = _RAND_211[255:0];
  _RAND_212 = {8{`RANDOM}};
  mem_212 = _RAND_212[255:0];
  _RAND_213 = {8{`RANDOM}};
  mem_213 = _RAND_213[255:0];
  _RAND_214 = {8{`RANDOM}};
  mem_214 = _RAND_214[255:0];
  _RAND_215 = {8{`RANDOM}};
  mem_215 = _RAND_215[255:0];
  _RAND_216 = {8{`RANDOM}};
  mem_216 = _RAND_216[255:0];
  _RAND_217 = {8{`RANDOM}};
  mem_217 = _RAND_217[255:0];
  _RAND_218 = {8{`RANDOM}};
  mem_218 = _RAND_218[255:0];
  _RAND_219 = {8{`RANDOM}};
  mem_219 = _RAND_219[255:0];
  _RAND_220 = {8{`RANDOM}};
  mem_220 = _RAND_220[255:0];
  _RAND_221 = {8{`RANDOM}};
  mem_221 = _RAND_221[255:0];
  _RAND_222 = {8{`RANDOM}};
  mem_222 = _RAND_222[255:0];
  _RAND_223 = {8{`RANDOM}};
  mem_223 = _RAND_223[255:0];
  _RAND_224 = {8{`RANDOM}};
  mem_224 = _RAND_224[255:0];
  _RAND_225 = {8{`RANDOM}};
  mem_225 = _RAND_225[255:0];
  _RAND_226 = {8{`RANDOM}};
  mem_226 = _RAND_226[255:0];
  _RAND_227 = {8{`RANDOM}};
  mem_227 = _RAND_227[255:0];
  _RAND_228 = {8{`RANDOM}};
  mem_228 = _RAND_228[255:0];
  _RAND_229 = {8{`RANDOM}};
  mem_229 = _RAND_229[255:0];
  _RAND_230 = {8{`RANDOM}};
  mem_230 = _RAND_230[255:0];
  _RAND_231 = {8{`RANDOM}};
  mem_231 = _RAND_231[255:0];
  _RAND_232 = {8{`RANDOM}};
  mem_232 = _RAND_232[255:0];
  _RAND_233 = {8{`RANDOM}};
  mem_233 = _RAND_233[255:0];
  _RAND_234 = {8{`RANDOM}};
  mem_234 = _RAND_234[255:0];
  _RAND_235 = {8{`RANDOM}};
  mem_235 = _RAND_235[255:0];
  _RAND_236 = {8{`RANDOM}};
  mem_236 = _RAND_236[255:0];
  _RAND_237 = {8{`RANDOM}};
  mem_237 = _RAND_237[255:0];
  _RAND_238 = {8{`RANDOM}};
  mem_238 = _RAND_238[255:0];
  _RAND_239 = {8{`RANDOM}};
  mem_239 = _RAND_239[255:0];
  _RAND_240 = {8{`RANDOM}};
  mem_240 = _RAND_240[255:0];
  _RAND_241 = {8{`RANDOM}};
  mem_241 = _RAND_241[255:0];
  _RAND_242 = {8{`RANDOM}};
  mem_242 = _RAND_242[255:0];
  _RAND_243 = {8{`RANDOM}};
  mem_243 = _RAND_243[255:0];
  _RAND_244 = {8{`RANDOM}};
  mem_244 = _RAND_244[255:0];
  _RAND_245 = {8{`RANDOM}};
  mem_245 = _RAND_245[255:0];
  _RAND_246 = {8{`RANDOM}};
  mem_246 = _RAND_246[255:0];
  _RAND_247 = {8{`RANDOM}};
  mem_247 = _RAND_247[255:0];
  _RAND_248 = {8{`RANDOM}};
  mem_248 = _RAND_248[255:0];
  _RAND_249 = {8{`RANDOM}};
  mem_249 = _RAND_249[255:0];
  _RAND_250 = {8{`RANDOM}};
  mem_250 = _RAND_250[255:0];
  _RAND_251 = {8{`RANDOM}};
  mem_251 = _RAND_251[255:0];
  _RAND_252 = {8{`RANDOM}};
  mem_252 = _RAND_252[255:0];
  _RAND_253 = {8{`RANDOM}};
  mem_253 = _RAND_253[255:0];
  _RAND_254 = {8{`RANDOM}};
  mem_254 = _RAND_254[255:0];
  _RAND_255 = {8{`RANDOM}};
  mem_255 = _RAND_255[255:0];
  _RAND_256 = {8{`RANDOM}};
  mem_256 = _RAND_256[255:0];
  _RAND_257 = {8{`RANDOM}};
  mem_257 = _RAND_257[255:0];
  _RAND_258 = {8{`RANDOM}};
  mem_258 = _RAND_258[255:0];
  _RAND_259 = {8{`RANDOM}};
  mem_259 = _RAND_259[255:0];
  _RAND_260 = {8{`RANDOM}};
  mem_260 = _RAND_260[255:0];
  _RAND_261 = {8{`RANDOM}};
  mem_261 = _RAND_261[255:0];
  _RAND_262 = {8{`RANDOM}};
  mem_262 = _RAND_262[255:0];
  _RAND_263 = {8{`RANDOM}};
  mem_263 = _RAND_263[255:0];
  _RAND_264 = {8{`RANDOM}};
  mem_264 = _RAND_264[255:0];
  _RAND_265 = {8{`RANDOM}};
  mem_265 = _RAND_265[255:0];
  _RAND_266 = {8{`RANDOM}};
  mem_266 = _RAND_266[255:0];
  _RAND_267 = {8{`RANDOM}};
  mem_267 = _RAND_267[255:0];
  _RAND_268 = {8{`RANDOM}};
  mem_268 = _RAND_268[255:0];
  _RAND_269 = {8{`RANDOM}};
  mem_269 = _RAND_269[255:0];
  _RAND_270 = {8{`RANDOM}};
  mem_270 = _RAND_270[255:0];
  _RAND_271 = {8{`RANDOM}};
  mem_271 = _RAND_271[255:0];
  _RAND_272 = {8{`RANDOM}};
  mem_272 = _RAND_272[255:0];
  _RAND_273 = {8{`RANDOM}};
  mem_273 = _RAND_273[255:0];
  _RAND_274 = {8{`RANDOM}};
  mem_274 = _RAND_274[255:0];
  _RAND_275 = {8{`RANDOM}};
  mem_275 = _RAND_275[255:0];
  _RAND_276 = {8{`RANDOM}};
  mem_276 = _RAND_276[255:0];
  _RAND_277 = {8{`RANDOM}};
  mem_277 = _RAND_277[255:0];
  _RAND_278 = {8{`RANDOM}};
  mem_278 = _RAND_278[255:0];
  _RAND_279 = {8{`RANDOM}};
  mem_279 = _RAND_279[255:0];
  _RAND_280 = {8{`RANDOM}};
  mem_280 = _RAND_280[255:0];
  _RAND_281 = {8{`RANDOM}};
  mem_281 = _RAND_281[255:0];
  _RAND_282 = {8{`RANDOM}};
  mem_282 = _RAND_282[255:0];
  _RAND_283 = {8{`RANDOM}};
  mem_283 = _RAND_283[255:0];
  _RAND_284 = {8{`RANDOM}};
  mem_284 = _RAND_284[255:0];
  _RAND_285 = {8{`RANDOM}};
  mem_285 = _RAND_285[255:0];
  _RAND_286 = {8{`RANDOM}};
  mem_286 = _RAND_286[255:0];
  _RAND_287 = {8{`RANDOM}};
  mem_287 = _RAND_287[255:0];
  _RAND_288 = {8{`RANDOM}};
  mem_288 = _RAND_288[255:0];
  _RAND_289 = {8{`RANDOM}};
  mem_289 = _RAND_289[255:0];
  _RAND_290 = {8{`RANDOM}};
  mem_290 = _RAND_290[255:0];
  _RAND_291 = {8{`RANDOM}};
  mem_291 = _RAND_291[255:0];
  _RAND_292 = {8{`RANDOM}};
  mem_292 = _RAND_292[255:0];
  _RAND_293 = {8{`RANDOM}};
  mem_293 = _RAND_293[255:0];
  _RAND_294 = {8{`RANDOM}};
  mem_294 = _RAND_294[255:0];
  _RAND_295 = {8{`RANDOM}};
  mem_295 = _RAND_295[255:0];
  _RAND_296 = {8{`RANDOM}};
  mem_296 = _RAND_296[255:0];
  _RAND_297 = {8{`RANDOM}};
  mem_297 = _RAND_297[255:0];
  _RAND_298 = {8{`RANDOM}};
  mem_298 = _RAND_298[255:0];
  _RAND_299 = {8{`RANDOM}};
  mem_299 = _RAND_299[255:0];
  _RAND_300 = {8{`RANDOM}};
  mem_300 = _RAND_300[255:0];
  _RAND_301 = {8{`RANDOM}};
  mem_301 = _RAND_301[255:0];
  _RAND_302 = {8{`RANDOM}};
  mem_302 = _RAND_302[255:0];
  _RAND_303 = {8{`RANDOM}};
  mem_303 = _RAND_303[255:0];
  _RAND_304 = {8{`RANDOM}};
  mem_304 = _RAND_304[255:0];
  _RAND_305 = {8{`RANDOM}};
  mem_305 = _RAND_305[255:0];
  _RAND_306 = {8{`RANDOM}};
  mem_306 = _RAND_306[255:0];
  _RAND_307 = {8{`RANDOM}};
  mem_307 = _RAND_307[255:0];
  _RAND_308 = {8{`RANDOM}};
  mem_308 = _RAND_308[255:0];
  _RAND_309 = {8{`RANDOM}};
  mem_309 = _RAND_309[255:0];
  _RAND_310 = {8{`RANDOM}};
  mem_310 = _RAND_310[255:0];
  _RAND_311 = {8{`RANDOM}};
  mem_311 = _RAND_311[255:0];
  _RAND_312 = {8{`RANDOM}};
  mem_312 = _RAND_312[255:0];
  _RAND_313 = {8{`RANDOM}};
  mem_313 = _RAND_313[255:0];
  _RAND_314 = {8{`RANDOM}};
  mem_314 = _RAND_314[255:0];
  _RAND_315 = {8{`RANDOM}};
  mem_315 = _RAND_315[255:0];
  _RAND_316 = {8{`RANDOM}};
  mem_316 = _RAND_316[255:0];
  _RAND_317 = {8{`RANDOM}};
  mem_317 = _RAND_317[255:0];
  _RAND_318 = {8{`RANDOM}};
  mem_318 = _RAND_318[255:0];
  _RAND_319 = {8{`RANDOM}};
  mem_319 = _RAND_319[255:0];
  _RAND_320 = {8{`RANDOM}};
  mem_320 = _RAND_320[255:0];
  _RAND_321 = {8{`RANDOM}};
  mem_321 = _RAND_321[255:0];
  _RAND_322 = {8{`RANDOM}};
  mem_322 = _RAND_322[255:0];
  _RAND_323 = {8{`RANDOM}};
  mem_323 = _RAND_323[255:0];
  _RAND_324 = {8{`RANDOM}};
  mem_324 = _RAND_324[255:0];
  _RAND_325 = {8{`RANDOM}};
  mem_325 = _RAND_325[255:0];
  _RAND_326 = {8{`RANDOM}};
  mem_326 = _RAND_326[255:0];
  _RAND_327 = {8{`RANDOM}};
  mem_327 = _RAND_327[255:0];
  _RAND_328 = {8{`RANDOM}};
  mem_328 = _RAND_328[255:0];
  _RAND_329 = {8{`RANDOM}};
  mem_329 = _RAND_329[255:0];
  _RAND_330 = {8{`RANDOM}};
  mem_330 = _RAND_330[255:0];
  _RAND_331 = {8{`RANDOM}};
  mem_331 = _RAND_331[255:0];
  _RAND_332 = {8{`RANDOM}};
  mem_332 = _RAND_332[255:0];
  _RAND_333 = {8{`RANDOM}};
  mem_333 = _RAND_333[255:0];
  _RAND_334 = {8{`RANDOM}};
  mem_334 = _RAND_334[255:0];
  _RAND_335 = {8{`RANDOM}};
  mem_335 = _RAND_335[255:0];
  _RAND_336 = {8{`RANDOM}};
  mem_336 = _RAND_336[255:0];
  _RAND_337 = {8{`RANDOM}};
  mem_337 = _RAND_337[255:0];
  _RAND_338 = {8{`RANDOM}};
  mem_338 = _RAND_338[255:0];
  _RAND_339 = {8{`RANDOM}};
  mem_339 = _RAND_339[255:0];
  _RAND_340 = {8{`RANDOM}};
  mem_340 = _RAND_340[255:0];
  _RAND_341 = {8{`RANDOM}};
  mem_341 = _RAND_341[255:0];
  _RAND_342 = {8{`RANDOM}};
  mem_342 = _RAND_342[255:0];
  _RAND_343 = {8{`RANDOM}};
  mem_343 = _RAND_343[255:0];
  _RAND_344 = {8{`RANDOM}};
  mem_344 = _RAND_344[255:0];
  _RAND_345 = {8{`RANDOM}};
  mem_345 = _RAND_345[255:0];
  _RAND_346 = {8{`RANDOM}};
  mem_346 = _RAND_346[255:0];
  _RAND_347 = {8{`RANDOM}};
  mem_347 = _RAND_347[255:0];
  _RAND_348 = {8{`RANDOM}};
  mem_348 = _RAND_348[255:0];
  _RAND_349 = {8{`RANDOM}};
  mem_349 = _RAND_349[255:0];
  _RAND_350 = {8{`RANDOM}};
  mem_350 = _RAND_350[255:0];
  _RAND_351 = {8{`RANDOM}};
  mem_351 = _RAND_351[255:0];
  _RAND_352 = {8{`RANDOM}};
  mem_352 = _RAND_352[255:0];
  _RAND_353 = {8{`RANDOM}};
  mem_353 = _RAND_353[255:0];
  _RAND_354 = {8{`RANDOM}};
  mem_354 = _RAND_354[255:0];
  _RAND_355 = {8{`RANDOM}};
  mem_355 = _RAND_355[255:0];
  _RAND_356 = {8{`RANDOM}};
  mem_356 = _RAND_356[255:0];
  _RAND_357 = {8{`RANDOM}};
  mem_357 = _RAND_357[255:0];
  _RAND_358 = {8{`RANDOM}};
  mem_358 = _RAND_358[255:0];
  _RAND_359 = {8{`RANDOM}};
  mem_359 = _RAND_359[255:0];
  _RAND_360 = {8{`RANDOM}};
  mem_360 = _RAND_360[255:0];
  _RAND_361 = {8{`RANDOM}};
  mem_361 = _RAND_361[255:0];
  _RAND_362 = {8{`RANDOM}};
  mem_362 = _RAND_362[255:0];
  _RAND_363 = {8{`RANDOM}};
  mem_363 = _RAND_363[255:0];
  _RAND_364 = {8{`RANDOM}};
  mem_364 = _RAND_364[255:0];
  _RAND_365 = {8{`RANDOM}};
  mem_365 = _RAND_365[255:0];
  _RAND_366 = {8{`RANDOM}};
  mem_366 = _RAND_366[255:0];
  _RAND_367 = {8{`RANDOM}};
  mem_367 = _RAND_367[255:0];
  _RAND_368 = {8{`RANDOM}};
  mem_368 = _RAND_368[255:0];
  _RAND_369 = {8{`RANDOM}};
  mem_369 = _RAND_369[255:0];
  _RAND_370 = {8{`RANDOM}};
  mem_370 = _RAND_370[255:0];
  _RAND_371 = {8{`RANDOM}};
  mem_371 = _RAND_371[255:0];
  _RAND_372 = {8{`RANDOM}};
  mem_372 = _RAND_372[255:0];
  _RAND_373 = {8{`RANDOM}};
  mem_373 = _RAND_373[255:0];
  _RAND_374 = {8{`RANDOM}};
  mem_374 = _RAND_374[255:0];
  _RAND_375 = {8{`RANDOM}};
  mem_375 = _RAND_375[255:0];
  _RAND_376 = {8{`RANDOM}};
  mem_376 = _RAND_376[255:0];
  _RAND_377 = {8{`RANDOM}};
  mem_377 = _RAND_377[255:0];
  _RAND_378 = {8{`RANDOM}};
  mem_378 = _RAND_378[255:0];
  _RAND_379 = {8{`RANDOM}};
  mem_379 = _RAND_379[255:0];
  _RAND_380 = {8{`RANDOM}};
  mem_380 = _RAND_380[255:0];
  _RAND_381 = {8{`RANDOM}};
  mem_381 = _RAND_381[255:0];
  _RAND_382 = {8{`RANDOM}};
  mem_382 = _RAND_382[255:0];
  _RAND_383 = {8{`RANDOM}};
  mem_383 = _RAND_383[255:0];
  _RAND_384 = {8{`RANDOM}};
  mem_384 = _RAND_384[255:0];
  _RAND_385 = {8{`RANDOM}};
  mem_385 = _RAND_385[255:0];
  _RAND_386 = {8{`RANDOM}};
  mem_386 = _RAND_386[255:0];
  _RAND_387 = {8{`RANDOM}};
  mem_387 = _RAND_387[255:0];
  _RAND_388 = {8{`RANDOM}};
  mem_388 = _RAND_388[255:0];
  _RAND_389 = {8{`RANDOM}};
  mem_389 = _RAND_389[255:0];
  _RAND_390 = {8{`RANDOM}};
  mem_390 = _RAND_390[255:0];
  _RAND_391 = {8{`RANDOM}};
  mem_391 = _RAND_391[255:0];
  _RAND_392 = {8{`RANDOM}};
  mem_392 = _RAND_392[255:0];
  _RAND_393 = {8{`RANDOM}};
  mem_393 = _RAND_393[255:0];
  _RAND_394 = {8{`RANDOM}};
  mem_394 = _RAND_394[255:0];
  _RAND_395 = {8{`RANDOM}};
  mem_395 = _RAND_395[255:0];
  _RAND_396 = {8{`RANDOM}};
  mem_396 = _RAND_396[255:0];
  _RAND_397 = {8{`RANDOM}};
  mem_397 = _RAND_397[255:0];
  _RAND_398 = {8{`RANDOM}};
  mem_398 = _RAND_398[255:0];
  _RAND_399 = {8{`RANDOM}};
  mem_399 = _RAND_399[255:0];
  _RAND_400 = {8{`RANDOM}};
  mem_400 = _RAND_400[255:0];
  _RAND_401 = {8{`RANDOM}};
  mem_401 = _RAND_401[255:0];
  _RAND_402 = {8{`RANDOM}};
  mem_402 = _RAND_402[255:0];
  _RAND_403 = {8{`RANDOM}};
  mem_403 = _RAND_403[255:0];
  _RAND_404 = {8{`RANDOM}};
  mem_404 = _RAND_404[255:0];
  _RAND_405 = {8{`RANDOM}};
  mem_405 = _RAND_405[255:0];
  _RAND_406 = {8{`RANDOM}};
  mem_406 = _RAND_406[255:0];
  _RAND_407 = {8{`RANDOM}};
  mem_407 = _RAND_407[255:0];
  _RAND_408 = {8{`RANDOM}};
  mem_408 = _RAND_408[255:0];
  _RAND_409 = {8{`RANDOM}};
  mem_409 = _RAND_409[255:0];
  _RAND_410 = {8{`RANDOM}};
  mem_410 = _RAND_410[255:0];
  _RAND_411 = {8{`RANDOM}};
  mem_411 = _RAND_411[255:0];
  _RAND_412 = {8{`RANDOM}};
  mem_412 = _RAND_412[255:0];
  _RAND_413 = {8{`RANDOM}};
  mem_413 = _RAND_413[255:0];
  _RAND_414 = {8{`RANDOM}};
  mem_414 = _RAND_414[255:0];
  _RAND_415 = {8{`RANDOM}};
  mem_415 = _RAND_415[255:0];
  _RAND_416 = {8{`RANDOM}};
  mem_416 = _RAND_416[255:0];
  _RAND_417 = {8{`RANDOM}};
  mem_417 = _RAND_417[255:0];
  _RAND_418 = {8{`RANDOM}};
  mem_418 = _RAND_418[255:0];
  _RAND_419 = {8{`RANDOM}};
  mem_419 = _RAND_419[255:0];
  _RAND_420 = {8{`RANDOM}};
  mem_420 = _RAND_420[255:0];
  _RAND_421 = {8{`RANDOM}};
  mem_421 = _RAND_421[255:0];
  _RAND_422 = {8{`RANDOM}};
  mem_422 = _RAND_422[255:0];
  _RAND_423 = {8{`RANDOM}};
  mem_423 = _RAND_423[255:0];
  _RAND_424 = {8{`RANDOM}};
  mem_424 = _RAND_424[255:0];
  _RAND_425 = {8{`RANDOM}};
  mem_425 = _RAND_425[255:0];
  _RAND_426 = {8{`RANDOM}};
  mem_426 = _RAND_426[255:0];
  _RAND_427 = {8{`RANDOM}};
  mem_427 = _RAND_427[255:0];
  _RAND_428 = {8{`RANDOM}};
  mem_428 = _RAND_428[255:0];
  _RAND_429 = {8{`RANDOM}};
  mem_429 = _RAND_429[255:0];
  _RAND_430 = {8{`RANDOM}};
  mem_430 = _RAND_430[255:0];
  _RAND_431 = {8{`RANDOM}};
  mem_431 = _RAND_431[255:0];
  _RAND_432 = {8{`RANDOM}};
  mem_432 = _RAND_432[255:0];
  _RAND_433 = {8{`RANDOM}};
  mem_433 = _RAND_433[255:0];
  _RAND_434 = {8{`RANDOM}};
  mem_434 = _RAND_434[255:0];
  _RAND_435 = {8{`RANDOM}};
  mem_435 = _RAND_435[255:0];
  _RAND_436 = {8{`RANDOM}};
  mem_436 = _RAND_436[255:0];
  _RAND_437 = {8{`RANDOM}};
  mem_437 = _RAND_437[255:0];
  _RAND_438 = {8{`RANDOM}};
  mem_438 = _RAND_438[255:0];
  _RAND_439 = {8{`RANDOM}};
  mem_439 = _RAND_439[255:0];
  _RAND_440 = {8{`RANDOM}};
  mem_440 = _RAND_440[255:0];
  _RAND_441 = {8{`RANDOM}};
  mem_441 = _RAND_441[255:0];
  _RAND_442 = {8{`RANDOM}};
  mem_442 = _RAND_442[255:0];
  _RAND_443 = {8{`RANDOM}};
  mem_443 = _RAND_443[255:0];
  _RAND_444 = {8{`RANDOM}};
  mem_444 = _RAND_444[255:0];
  _RAND_445 = {8{`RANDOM}};
  mem_445 = _RAND_445[255:0];
  _RAND_446 = {8{`RANDOM}};
  mem_446 = _RAND_446[255:0];
  _RAND_447 = {8{`RANDOM}};
  mem_447 = _RAND_447[255:0];
  _RAND_448 = {8{`RANDOM}};
  mem_448 = _RAND_448[255:0];
  _RAND_449 = {8{`RANDOM}};
  mem_449 = _RAND_449[255:0];
  _RAND_450 = {8{`RANDOM}};
  mem_450 = _RAND_450[255:0];
  _RAND_451 = {8{`RANDOM}};
  mem_451 = _RAND_451[255:0];
  _RAND_452 = {8{`RANDOM}};
  mem_452 = _RAND_452[255:0];
  _RAND_453 = {8{`RANDOM}};
  mem_453 = _RAND_453[255:0];
  _RAND_454 = {8{`RANDOM}};
  mem_454 = _RAND_454[255:0];
  _RAND_455 = {8{`RANDOM}};
  mem_455 = _RAND_455[255:0];
  _RAND_456 = {8{`RANDOM}};
  mem_456 = _RAND_456[255:0];
  _RAND_457 = {8{`RANDOM}};
  mem_457 = _RAND_457[255:0];
  _RAND_458 = {8{`RANDOM}};
  mem_458 = _RAND_458[255:0];
  _RAND_459 = {8{`RANDOM}};
  mem_459 = _RAND_459[255:0];
  _RAND_460 = {8{`RANDOM}};
  mem_460 = _RAND_460[255:0];
  _RAND_461 = {8{`RANDOM}};
  mem_461 = _RAND_461[255:0];
  _RAND_462 = {8{`RANDOM}};
  mem_462 = _RAND_462[255:0];
  _RAND_463 = {8{`RANDOM}};
  mem_463 = _RAND_463[255:0];
  _RAND_464 = {8{`RANDOM}};
  mem_464 = _RAND_464[255:0];
  _RAND_465 = {8{`RANDOM}};
  mem_465 = _RAND_465[255:0];
  _RAND_466 = {8{`RANDOM}};
  mem_466 = _RAND_466[255:0];
  _RAND_467 = {8{`RANDOM}};
  mem_467 = _RAND_467[255:0];
  _RAND_468 = {8{`RANDOM}};
  mem_468 = _RAND_468[255:0];
  _RAND_469 = {8{`RANDOM}};
  mem_469 = _RAND_469[255:0];
  _RAND_470 = {8{`RANDOM}};
  mem_470 = _RAND_470[255:0];
  _RAND_471 = {8{`RANDOM}};
  mem_471 = _RAND_471[255:0];
  _RAND_472 = {8{`RANDOM}};
  mem_472 = _RAND_472[255:0];
  _RAND_473 = {8{`RANDOM}};
  mem_473 = _RAND_473[255:0];
  _RAND_474 = {8{`RANDOM}};
  mem_474 = _RAND_474[255:0];
  _RAND_475 = {8{`RANDOM}};
  mem_475 = _RAND_475[255:0];
  _RAND_476 = {8{`RANDOM}};
  mem_476 = _RAND_476[255:0];
  _RAND_477 = {8{`RANDOM}};
  mem_477 = _RAND_477[255:0];
  _RAND_478 = {8{`RANDOM}};
  mem_478 = _RAND_478[255:0];
  _RAND_479 = {8{`RANDOM}};
  mem_479 = _RAND_479[255:0];
  _RAND_480 = {8{`RANDOM}};
  mem_480 = _RAND_480[255:0];
  _RAND_481 = {8{`RANDOM}};
  mem_481 = _RAND_481[255:0];
  _RAND_482 = {8{`RANDOM}};
  mem_482 = _RAND_482[255:0];
  _RAND_483 = {8{`RANDOM}};
  mem_483 = _RAND_483[255:0];
  _RAND_484 = {8{`RANDOM}};
  mem_484 = _RAND_484[255:0];
  _RAND_485 = {8{`RANDOM}};
  mem_485 = _RAND_485[255:0];
  _RAND_486 = {8{`RANDOM}};
  mem_486 = _RAND_486[255:0];
  _RAND_487 = {8{`RANDOM}};
  mem_487 = _RAND_487[255:0];
  _RAND_488 = {8{`RANDOM}};
  mem_488 = _RAND_488[255:0];
  _RAND_489 = {8{`RANDOM}};
  mem_489 = _RAND_489[255:0];
  _RAND_490 = {8{`RANDOM}};
  mem_490 = _RAND_490[255:0];
  _RAND_491 = {8{`RANDOM}};
  mem_491 = _RAND_491[255:0];
  _RAND_492 = {8{`RANDOM}};
  mem_492 = _RAND_492[255:0];
  _RAND_493 = {8{`RANDOM}};
  mem_493 = _RAND_493[255:0];
  _RAND_494 = {8{`RANDOM}};
  mem_494 = _RAND_494[255:0];
  _RAND_495 = {8{`RANDOM}};
  mem_495 = _RAND_495[255:0];
  _RAND_496 = {8{`RANDOM}};
  mem_496 = _RAND_496[255:0];
  _RAND_497 = {8{`RANDOM}};
  mem_497 = _RAND_497[255:0];
  _RAND_498 = {8{`RANDOM}};
  mem_498 = _RAND_498[255:0];
  _RAND_499 = {8{`RANDOM}};
  mem_499 = _RAND_499[255:0];
  _RAND_500 = {8{`RANDOM}};
  mem_500 = _RAND_500[255:0];
  _RAND_501 = {8{`RANDOM}};
  mem_501 = _RAND_501[255:0];
  _RAND_502 = {8{`RANDOM}};
  mem_502 = _RAND_502[255:0];
  _RAND_503 = {8{`RANDOM}};
  mem_503 = _RAND_503[255:0];
  _RAND_504 = {8{`RANDOM}};
  mem_504 = _RAND_504[255:0];
  _RAND_505 = {8{`RANDOM}};
  mem_505 = _RAND_505[255:0];
  _RAND_506 = {8{`RANDOM}};
  mem_506 = _RAND_506[255:0];
  _RAND_507 = {8{`RANDOM}};
  mem_507 = _RAND_507[255:0];
  _RAND_508 = {8{`RANDOM}};
  mem_508 = _RAND_508[255:0];
  _RAND_509 = {8{`RANDOM}};
  mem_509 = _RAND_509[255:0];
  _RAND_510 = {8{`RANDOM}};
  mem_510 = _RAND_510[255:0];
  _RAND_511 = {8{`RANDOM}};
  mem_511 = _RAND_511[255:0];
  _RAND_512 = {8{`RANDOM}};
  io_dout_REG = _RAND_512[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinglePortBRAM(
  input          clock,
  input          reset,
  input          io_we,
  input  [8:0]   io_addr,
  input  [255:0] io_din,
  output [255:0] io_dout
);
  wire  sim_single_port_bram_clock; // @[RAMWrapper.scala 275:38]
  wire  sim_single_port_bram_reset; // @[RAMWrapper.scala 275:38]
  wire  sim_single_port_bram_io_we; // @[RAMWrapper.scala 275:38]
  wire [8:0] sim_single_port_bram_io_addr; // @[RAMWrapper.scala 275:38]
  wire [255:0] sim_single_port_bram_io_din; // @[RAMWrapper.scala 275:38]
  wire [255:0] sim_single_port_bram_io_dout; // @[RAMWrapper.scala 275:38]
  SimSinglePortBRAM sim_single_port_bram ( // @[RAMWrapper.scala 275:38]
    .clock(sim_single_port_bram_clock),
    .reset(sim_single_port_bram_reset),
    .io_we(sim_single_port_bram_io_we),
    .io_addr(sim_single_port_bram_io_addr),
    .io_din(sim_single_port_bram_io_din),
    .io_dout(sim_single_port_bram_io_dout)
  );
  assign io_dout = sim_single_port_bram_io_dout; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_clock = clock;
  assign sim_single_port_bram_reset = reset;
  assign sim_single_port_bram_io_we = io_we; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_io_addr = io_addr; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_io_din = io_din; // @[RAMWrapper.scala 276:29]
endmodule
module SimSinglePortBRAM_1(
  input         clock,
  input         reset,
  input         io_we,
  input  [8:0]  io_addr,
  input  [18:0] io_din,
  output [18:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] mem_0; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_1; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_2; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_3; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_4; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_5; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_6; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_7; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_8; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_9; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_10; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_11; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_12; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_13; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_14; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_15; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_16; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_17; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_18; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_19; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_20; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_21; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_22; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_23; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_24; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_25; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_26; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_27; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_28; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_29; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_30; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_31; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_32; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_33; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_34; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_35; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_36; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_37; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_38; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_39; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_40; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_41; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_42; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_43; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_44; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_45; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_46; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_47; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_48; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_49; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_50; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_51; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_52; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_53; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_54; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_55; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_56; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_57; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_58; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_59; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_60; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_61; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_62; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_63; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_64; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_65; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_66; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_67; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_68; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_69; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_70; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_71; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_72; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_73; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_74; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_75; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_76; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_77; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_78; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_79; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_80; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_81; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_82; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_83; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_84; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_85; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_86; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_87; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_88; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_89; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_90; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_91; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_92; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_93; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_94; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_95; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_96; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_97; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_98; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_99; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_100; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_101; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_102; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_103; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_104; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_105; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_106; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_107; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_108; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_109; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_110; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_111; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_112; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_113; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_114; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_115; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_116; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_117; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_118; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_119; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_120; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_121; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_122; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_123; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_124; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_125; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_126; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_127; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_128; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_129; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_130; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_131; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_132; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_133; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_134; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_135; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_136; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_137; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_138; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_139; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_140; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_141; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_142; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_143; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_144; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_145; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_146; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_147; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_148; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_149; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_150; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_151; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_152; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_153; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_154; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_155; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_156; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_157; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_158; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_159; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_160; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_161; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_162; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_163; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_164; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_165; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_166; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_167; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_168; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_169; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_170; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_171; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_172; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_173; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_174; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_175; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_176; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_177; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_178; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_179; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_180; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_181; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_182; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_183; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_184; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_185; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_186; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_187; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_188; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_189; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_190; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_191; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_192; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_193; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_194; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_195; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_196; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_197; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_198; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_199; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_200; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_201; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_202; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_203; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_204; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_205; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_206; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_207; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_208; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_209; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_210; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_211; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_212; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_213; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_214; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_215; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_216; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_217; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_218; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_219; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_220; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_221; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_222; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_223; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_224; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_225; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_226; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_227; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_228; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_229; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_230; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_231; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_232; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_233; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_234; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_235; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_236; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_237; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_238; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_239; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_240; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_241; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_242; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_243; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_244; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_245; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_246; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_247; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_248; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_249; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_250; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_251; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_252; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_253; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_254; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_255; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_256; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_257; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_258; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_259; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_260; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_261; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_262; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_263; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_264; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_265; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_266; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_267; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_268; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_269; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_270; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_271; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_272; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_273; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_274; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_275; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_276; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_277; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_278; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_279; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_280; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_281; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_282; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_283; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_284; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_285; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_286; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_287; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_288; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_289; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_290; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_291; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_292; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_293; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_294; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_295; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_296; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_297; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_298; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_299; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_300; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_301; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_302; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_303; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_304; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_305; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_306; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_307; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_308; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_309; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_310; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_311; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_312; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_313; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_314; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_315; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_316; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_317; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_318; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_319; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_320; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_321; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_322; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_323; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_324; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_325; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_326; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_327; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_328; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_329; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_330; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_331; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_332; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_333; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_334; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_335; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_336; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_337; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_338; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_339; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_340; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_341; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_342; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_343; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_344; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_345; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_346; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_347; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_348; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_349; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_350; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_351; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_352; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_353; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_354; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_355; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_356; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_357; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_358; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_359; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_360; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_361; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_362; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_363; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_364; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_365; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_366; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_367; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_368; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_369; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_370; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_371; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_372; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_373; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_374; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_375; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_376; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_377; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_378; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_379; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_380; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_381; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_382; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_383; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_384; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_385; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_386; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_387; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_388; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_389; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_390; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_391; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_392; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_393; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_394; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_395; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_396; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_397; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_398; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_399; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_400; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_401; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_402; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_403; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_404; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_405; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_406; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_407; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_408; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_409; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_410; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_411; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_412; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_413; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_414; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_415; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_416; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_417; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_418; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_419; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_420; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_421; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_422; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_423; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_424; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_425; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_426; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_427; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_428; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_429; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_430; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_431; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_432; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_433; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_434; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_435; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_436; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_437; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_438; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_439; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_440; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_441; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_442; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_443; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_444; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_445; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_446; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_447; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_448; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_449; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_450; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_451; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_452; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_453; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_454; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_455; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_456; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_457; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_458; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_459; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_460; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_461; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_462; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_463; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_464; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_465; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_466; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_467; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_468; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_469; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_470; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_471; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_472; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_473; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_474; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_475; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_476; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_477; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_478; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_479; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_480; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_481; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_482; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_483; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_484; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_485; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_486; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_487; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_488; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_489; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_490; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_491; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_492; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_493; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_494; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_495; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_496; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_497; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_498; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_499; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_500; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_501; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_502; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_503; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_504; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_505; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_506; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_507; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_508; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_509; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_510; // @[RAMWrapper.scala 286:20]
  reg [18:0] mem_511; // @[RAMWrapper.scala 286:20]
  reg [18:0] io_dout_REG; // @[RAMWrapper.scala 288:21]
  wire [18:0] _GEN_1 = 9'h1 == io_addr ? mem_1 : mem_0; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_2 = 9'h2 == io_addr ? mem_2 : _GEN_1; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_3 = 9'h3 == io_addr ? mem_3 : _GEN_2; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_4 = 9'h4 == io_addr ? mem_4 : _GEN_3; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_5 = 9'h5 == io_addr ? mem_5 : _GEN_4; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_6 = 9'h6 == io_addr ? mem_6 : _GEN_5; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_7 = 9'h7 == io_addr ? mem_7 : _GEN_6; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_8 = 9'h8 == io_addr ? mem_8 : _GEN_7; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_9 = 9'h9 == io_addr ? mem_9 : _GEN_8; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_10 = 9'ha == io_addr ? mem_10 : _GEN_9; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_11 = 9'hb == io_addr ? mem_11 : _GEN_10; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_12 = 9'hc == io_addr ? mem_12 : _GEN_11; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_13 = 9'hd == io_addr ? mem_13 : _GEN_12; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_14 = 9'he == io_addr ? mem_14 : _GEN_13; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_15 = 9'hf == io_addr ? mem_15 : _GEN_14; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_16 = 9'h10 == io_addr ? mem_16 : _GEN_15; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_17 = 9'h11 == io_addr ? mem_17 : _GEN_16; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_18 = 9'h12 == io_addr ? mem_18 : _GEN_17; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_19 = 9'h13 == io_addr ? mem_19 : _GEN_18; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_20 = 9'h14 == io_addr ? mem_20 : _GEN_19; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_21 = 9'h15 == io_addr ? mem_21 : _GEN_20; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_22 = 9'h16 == io_addr ? mem_22 : _GEN_21; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_23 = 9'h17 == io_addr ? mem_23 : _GEN_22; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_24 = 9'h18 == io_addr ? mem_24 : _GEN_23; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_25 = 9'h19 == io_addr ? mem_25 : _GEN_24; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_26 = 9'h1a == io_addr ? mem_26 : _GEN_25; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_27 = 9'h1b == io_addr ? mem_27 : _GEN_26; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_28 = 9'h1c == io_addr ? mem_28 : _GEN_27; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_29 = 9'h1d == io_addr ? mem_29 : _GEN_28; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_30 = 9'h1e == io_addr ? mem_30 : _GEN_29; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_31 = 9'h1f == io_addr ? mem_31 : _GEN_30; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_32 = 9'h20 == io_addr ? mem_32 : _GEN_31; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_33 = 9'h21 == io_addr ? mem_33 : _GEN_32; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_34 = 9'h22 == io_addr ? mem_34 : _GEN_33; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_35 = 9'h23 == io_addr ? mem_35 : _GEN_34; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_36 = 9'h24 == io_addr ? mem_36 : _GEN_35; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_37 = 9'h25 == io_addr ? mem_37 : _GEN_36; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_38 = 9'h26 == io_addr ? mem_38 : _GEN_37; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_39 = 9'h27 == io_addr ? mem_39 : _GEN_38; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_40 = 9'h28 == io_addr ? mem_40 : _GEN_39; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_41 = 9'h29 == io_addr ? mem_41 : _GEN_40; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_42 = 9'h2a == io_addr ? mem_42 : _GEN_41; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_43 = 9'h2b == io_addr ? mem_43 : _GEN_42; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_44 = 9'h2c == io_addr ? mem_44 : _GEN_43; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_45 = 9'h2d == io_addr ? mem_45 : _GEN_44; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_46 = 9'h2e == io_addr ? mem_46 : _GEN_45; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_47 = 9'h2f == io_addr ? mem_47 : _GEN_46; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_48 = 9'h30 == io_addr ? mem_48 : _GEN_47; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_49 = 9'h31 == io_addr ? mem_49 : _GEN_48; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_50 = 9'h32 == io_addr ? mem_50 : _GEN_49; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_51 = 9'h33 == io_addr ? mem_51 : _GEN_50; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_52 = 9'h34 == io_addr ? mem_52 : _GEN_51; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_53 = 9'h35 == io_addr ? mem_53 : _GEN_52; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_54 = 9'h36 == io_addr ? mem_54 : _GEN_53; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_55 = 9'h37 == io_addr ? mem_55 : _GEN_54; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_56 = 9'h38 == io_addr ? mem_56 : _GEN_55; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_57 = 9'h39 == io_addr ? mem_57 : _GEN_56; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_58 = 9'h3a == io_addr ? mem_58 : _GEN_57; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_59 = 9'h3b == io_addr ? mem_59 : _GEN_58; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_60 = 9'h3c == io_addr ? mem_60 : _GEN_59; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_61 = 9'h3d == io_addr ? mem_61 : _GEN_60; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_62 = 9'h3e == io_addr ? mem_62 : _GEN_61; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_63 = 9'h3f == io_addr ? mem_63 : _GEN_62; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_64 = 9'h40 == io_addr ? mem_64 : _GEN_63; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_65 = 9'h41 == io_addr ? mem_65 : _GEN_64; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_66 = 9'h42 == io_addr ? mem_66 : _GEN_65; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_67 = 9'h43 == io_addr ? mem_67 : _GEN_66; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_68 = 9'h44 == io_addr ? mem_68 : _GEN_67; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_69 = 9'h45 == io_addr ? mem_69 : _GEN_68; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_70 = 9'h46 == io_addr ? mem_70 : _GEN_69; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_71 = 9'h47 == io_addr ? mem_71 : _GEN_70; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_72 = 9'h48 == io_addr ? mem_72 : _GEN_71; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_73 = 9'h49 == io_addr ? mem_73 : _GEN_72; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_74 = 9'h4a == io_addr ? mem_74 : _GEN_73; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_75 = 9'h4b == io_addr ? mem_75 : _GEN_74; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_76 = 9'h4c == io_addr ? mem_76 : _GEN_75; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_77 = 9'h4d == io_addr ? mem_77 : _GEN_76; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_78 = 9'h4e == io_addr ? mem_78 : _GEN_77; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_79 = 9'h4f == io_addr ? mem_79 : _GEN_78; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_80 = 9'h50 == io_addr ? mem_80 : _GEN_79; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_81 = 9'h51 == io_addr ? mem_81 : _GEN_80; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_82 = 9'h52 == io_addr ? mem_82 : _GEN_81; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_83 = 9'h53 == io_addr ? mem_83 : _GEN_82; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_84 = 9'h54 == io_addr ? mem_84 : _GEN_83; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_85 = 9'h55 == io_addr ? mem_85 : _GEN_84; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_86 = 9'h56 == io_addr ? mem_86 : _GEN_85; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_87 = 9'h57 == io_addr ? mem_87 : _GEN_86; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_88 = 9'h58 == io_addr ? mem_88 : _GEN_87; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_89 = 9'h59 == io_addr ? mem_89 : _GEN_88; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_90 = 9'h5a == io_addr ? mem_90 : _GEN_89; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_91 = 9'h5b == io_addr ? mem_91 : _GEN_90; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_92 = 9'h5c == io_addr ? mem_92 : _GEN_91; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_93 = 9'h5d == io_addr ? mem_93 : _GEN_92; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_94 = 9'h5e == io_addr ? mem_94 : _GEN_93; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_95 = 9'h5f == io_addr ? mem_95 : _GEN_94; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_96 = 9'h60 == io_addr ? mem_96 : _GEN_95; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_97 = 9'h61 == io_addr ? mem_97 : _GEN_96; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_98 = 9'h62 == io_addr ? mem_98 : _GEN_97; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_99 = 9'h63 == io_addr ? mem_99 : _GEN_98; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_100 = 9'h64 == io_addr ? mem_100 : _GEN_99; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_101 = 9'h65 == io_addr ? mem_101 : _GEN_100; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_102 = 9'h66 == io_addr ? mem_102 : _GEN_101; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_103 = 9'h67 == io_addr ? mem_103 : _GEN_102; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_104 = 9'h68 == io_addr ? mem_104 : _GEN_103; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_105 = 9'h69 == io_addr ? mem_105 : _GEN_104; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_106 = 9'h6a == io_addr ? mem_106 : _GEN_105; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_107 = 9'h6b == io_addr ? mem_107 : _GEN_106; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_108 = 9'h6c == io_addr ? mem_108 : _GEN_107; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_109 = 9'h6d == io_addr ? mem_109 : _GEN_108; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_110 = 9'h6e == io_addr ? mem_110 : _GEN_109; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_111 = 9'h6f == io_addr ? mem_111 : _GEN_110; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_112 = 9'h70 == io_addr ? mem_112 : _GEN_111; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_113 = 9'h71 == io_addr ? mem_113 : _GEN_112; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_114 = 9'h72 == io_addr ? mem_114 : _GEN_113; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_115 = 9'h73 == io_addr ? mem_115 : _GEN_114; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_116 = 9'h74 == io_addr ? mem_116 : _GEN_115; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_117 = 9'h75 == io_addr ? mem_117 : _GEN_116; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_118 = 9'h76 == io_addr ? mem_118 : _GEN_117; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_119 = 9'h77 == io_addr ? mem_119 : _GEN_118; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_120 = 9'h78 == io_addr ? mem_120 : _GEN_119; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_121 = 9'h79 == io_addr ? mem_121 : _GEN_120; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_122 = 9'h7a == io_addr ? mem_122 : _GEN_121; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_123 = 9'h7b == io_addr ? mem_123 : _GEN_122; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_124 = 9'h7c == io_addr ? mem_124 : _GEN_123; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_125 = 9'h7d == io_addr ? mem_125 : _GEN_124; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_126 = 9'h7e == io_addr ? mem_126 : _GEN_125; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_127 = 9'h7f == io_addr ? mem_127 : _GEN_126; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_128 = 9'h80 == io_addr ? mem_128 : _GEN_127; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_129 = 9'h81 == io_addr ? mem_129 : _GEN_128; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_130 = 9'h82 == io_addr ? mem_130 : _GEN_129; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_131 = 9'h83 == io_addr ? mem_131 : _GEN_130; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_132 = 9'h84 == io_addr ? mem_132 : _GEN_131; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_133 = 9'h85 == io_addr ? mem_133 : _GEN_132; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_134 = 9'h86 == io_addr ? mem_134 : _GEN_133; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_135 = 9'h87 == io_addr ? mem_135 : _GEN_134; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_136 = 9'h88 == io_addr ? mem_136 : _GEN_135; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_137 = 9'h89 == io_addr ? mem_137 : _GEN_136; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_138 = 9'h8a == io_addr ? mem_138 : _GEN_137; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_139 = 9'h8b == io_addr ? mem_139 : _GEN_138; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_140 = 9'h8c == io_addr ? mem_140 : _GEN_139; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_141 = 9'h8d == io_addr ? mem_141 : _GEN_140; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_142 = 9'h8e == io_addr ? mem_142 : _GEN_141; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_143 = 9'h8f == io_addr ? mem_143 : _GEN_142; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_144 = 9'h90 == io_addr ? mem_144 : _GEN_143; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_145 = 9'h91 == io_addr ? mem_145 : _GEN_144; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_146 = 9'h92 == io_addr ? mem_146 : _GEN_145; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_147 = 9'h93 == io_addr ? mem_147 : _GEN_146; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_148 = 9'h94 == io_addr ? mem_148 : _GEN_147; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_149 = 9'h95 == io_addr ? mem_149 : _GEN_148; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_150 = 9'h96 == io_addr ? mem_150 : _GEN_149; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_151 = 9'h97 == io_addr ? mem_151 : _GEN_150; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_152 = 9'h98 == io_addr ? mem_152 : _GEN_151; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_153 = 9'h99 == io_addr ? mem_153 : _GEN_152; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_154 = 9'h9a == io_addr ? mem_154 : _GEN_153; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_155 = 9'h9b == io_addr ? mem_155 : _GEN_154; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_156 = 9'h9c == io_addr ? mem_156 : _GEN_155; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_157 = 9'h9d == io_addr ? mem_157 : _GEN_156; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_158 = 9'h9e == io_addr ? mem_158 : _GEN_157; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_159 = 9'h9f == io_addr ? mem_159 : _GEN_158; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_160 = 9'ha0 == io_addr ? mem_160 : _GEN_159; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_161 = 9'ha1 == io_addr ? mem_161 : _GEN_160; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_162 = 9'ha2 == io_addr ? mem_162 : _GEN_161; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_163 = 9'ha3 == io_addr ? mem_163 : _GEN_162; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_164 = 9'ha4 == io_addr ? mem_164 : _GEN_163; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_165 = 9'ha5 == io_addr ? mem_165 : _GEN_164; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_166 = 9'ha6 == io_addr ? mem_166 : _GEN_165; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_167 = 9'ha7 == io_addr ? mem_167 : _GEN_166; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_168 = 9'ha8 == io_addr ? mem_168 : _GEN_167; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_169 = 9'ha9 == io_addr ? mem_169 : _GEN_168; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_170 = 9'haa == io_addr ? mem_170 : _GEN_169; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_171 = 9'hab == io_addr ? mem_171 : _GEN_170; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_172 = 9'hac == io_addr ? mem_172 : _GEN_171; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_173 = 9'had == io_addr ? mem_173 : _GEN_172; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_174 = 9'hae == io_addr ? mem_174 : _GEN_173; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_175 = 9'haf == io_addr ? mem_175 : _GEN_174; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_176 = 9'hb0 == io_addr ? mem_176 : _GEN_175; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_177 = 9'hb1 == io_addr ? mem_177 : _GEN_176; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_178 = 9'hb2 == io_addr ? mem_178 : _GEN_177; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_179 = 9'hb3 == io_addr ? mem_179 : _GEN_178; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_180 = 9'hb4 == io_addr ? mem_180 : _GEN_179; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_181 = 9'hb5 == io_addr ? mem_181 : _GEN_180; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_182 = 9'hb6 == io_addr ? mem_182 : _GEN_181; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_183 = 9'hb7 == io_addr ? mem_183 : _GEN_182; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_184 = 9'hb8 == io_addr ? mem_184 : _GEN_183; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_185 = 9'hb9 == io_addr ? mem_185 : _GEN_184; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_186 = 9'hba == io_addr ? mem_186 : _GEN_185; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_187 = 9'hbb == io_addr ? mem_187 : _GEN_186; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_188 = 9'hbc == io_addr ? mem_188 : _GEN_187; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_189 = 9'hbd == io_addr ? mem_189 : _GEN_188; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_190 = 9'hbe == io_addr ? mem_190 : _GEN_189; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_191 = 9'hbf == io_addr ? mem_191 : _GEN_190; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_192 = 9'hc0 == io_addr ? mem_192 : _GEN_191; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_193 = 9'hc1 == io_addr ? mem_193 : _GEN_192; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_194 = 9'hc2 == io_addr ? mem_194 : _GEN_193; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_195 = 9'hc3 == io_addr ? mem_195 : _GEN_194; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_196 = 9'hc4 == io_addr ? mem_196 : _GEN_195; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_197 = 9'hc5 == io_addr ? mem_197 : _GEN_196; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_198 = 9'hc6 == io_addr ? mem_198 : _GEN_197; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_199 = 9'hc7 == io_addr ? mem_199 : _GEN_198; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_200 = 9'hc8 == io_addr ? mem_200 : _GEN_199; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_201 = 9'hc9 == io_addr ? mem_201 : _GEN_200; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_202 = 9'hca == io_addr ? mem_202 : _GEN_201; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_203 = 9'hcb == io_addr ? mem_203 : _GEN_202; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_204 = 9'hcc == io_addr ? mem_204 : _GEN_203; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_205 = 9'hcd == io_addr ? mem_205 : _GEN_204; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_206 = 9'hce == io_addr ? mem_206 : _GEN_205; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_207 = 9'hcf == io_addr ? mem_207 : _GEN_206; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_208 = 9'hd0 == io_addr ? mem_208 : _GEN_207; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_209 = 9'hd1 == io_addr ? mem_209 : _GEN_208; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_210 = 9'hd2 == io_addr ? mem_210 : _GEN_209; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_211 = 9'hd3 == io_addr ? mem_211 : _GEN_210; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_212 = 9'hd4 == io_addr ? mem_212 : _GEN_211; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_213 = 9'hd5 == io_addr ? mem_213 : _GEN_212; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_214 = 9'hd6 == io_addr ? mem_214 : _GEN_213; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_215 = 9'hd7 == io_addr ? mem_215 : _GEN_214; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_216 = 9'hd8 == io_addr ? mem_216 : _GEN_215; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_217 = 9'hd9 == io_addr ? mem_217 : _GEN_216; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_218 = 9'hda == io_addr ? mem_218 : _GEN_217; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_219 = 9'hdb == io_addr ? mem_219 : _GEN_218; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_220 = 9'hdc == io_addr ? mem_220 : _GEN_219; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_221 = 9'hdd == io_addr ? mem_221 : _GEN_220; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_222 = 9'hde == io_addr ? mem_222 : _GEN_221; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_223 = 9'hdf == io_addr ? mem_223 : _GEN_222; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_224 = 9'he0 == io_addr ? mem_224 : _GEN_223; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_225 = 9'he1 == io_addr ? mem_225 : _GEN_224; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_226 = 9'he2 == io_addr ? mem_226 : _GEN_225; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_227 = 9'he3 == io_addr ? mem_227 : _GEN_226; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_228 = 9'he4 == io_addr ? mem_228 : _GEN_227; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_229 = 9'he5 == io_addr ? mem_229 : _GEN_228; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_230 = 9'he6 == io_addr ? mem_230 : _GEN_229; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_231 = 9'he7 == io_addr ? mem_231 : _GEN_230; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_232 = 9'he8 == io_addr ? mem_232 : _GEN_231; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_233 = 9'he9 == io_addr ? mem_233 : _GEN_232; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_234 = 9'hea == io_addr ? mem_234 : _GEN_233; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_235 = 9'heb == io_addr ? mem_235 : _GEN_234; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_236 = 9'hec == io_addr ? mem_236 : _GEN_235; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_237 = 9'hed == io_addr ? mem_237 : _GEN_236; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_238 = 9'hee == io_addr ? mem_238 : _GEN_237; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_239 = 9'hef == io_addr ? mem_239 : _GEN_238; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_240 = 9'hf0 == io_addr ? mem_240 : _GEN_239; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_241 = 9'hf1 == io_addr ? mem_241 : _GEN_240; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_242 = 9'hf2 == io_addr ? mem_242 : _GEN_241; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_243 = 9'hf3 == io_addr ? mem_243 : _GEN_242; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_244 = 9'hf4 == io_addr ? mem_244 : _GEN_243; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_245 = 9'hf5 == io_addr ? mem_245 : _GEN_244; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_246 = 9'hf6 == io_addr ? mem_246 : _GEN_245; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_247 = 9'hf7 == io_addr ? mem_247 : _GEN_246; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_248 = 9'hf8 == io_addr ? mem_248 : _GEN_247; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_249 = 9'hf9 == io_addr ? mem_249 : _GEN_248; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_250 = 9'hfa == io_addr ? mem_250 : _GEN_249; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_251 = 9'hfb == io_addr ? mem_251 : _GEN_250; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_252 = 9'hfc == io_addr ? mem_252 : _GEN_251; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_253 = 9'hfd == io_addr ? mem_253 : _GEN_252; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_254 = 9'hfe == io_addr ? mem_254 : _GEN_253; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_255 = 9'hff == io_addr ? mem_255 : _GEN_254; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_256 = 9'h100 == io_addr ? mem_256 : _GEN_255; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_257 = 9'h101 == io_addr ? mem_257 : _GEN_256; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_258 = 9'h102 == io_addr ? mem_258 : _GEN_257; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_259 = 9'h103 == io_addr ? mem_259 : _GEN_258; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_260 = 9'h104 == io_addr ? mem_260 : _GEN_259; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_261 = 9'h105 == io_addr ? mem_261 : _GEN_260; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_262 = 9'h106 == io_addr ? mem_262 : _GEN_261; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_263 = 9'h107 == io_addr ? mem_263 : _GEN_262; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_264 = 9'h108 == io_addr ? mem_264 : _GEN_263; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_265 = 9'h109 == io_addr ? mem_265 : _GEN_264; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_266 = 9'h10a == io_addr ? mem_266 : _GEN_265; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_267 = 9'h10b == io_addr ? mem_267 : _GEN_266; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_268 = 9'h10c == io_addr ? mem_268 : _GEN_267; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_269 = 9'h10d == io_addr ? mem_269 : _GEN_268; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_270 = 9'h10e == io_addr ? mem_270 : _GEN_269; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_271 = 9'h10f == io_addr ? mem_271 : _GEN_270; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_272 = 9'h110 == io_addr ? mem_272 : _GEN_271; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_273 = 9'h111 == io_addr ? mem_273 : _GEN_272; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_274 = 9'h112 == io_addr ? mem_274 : _GEN_273; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_275 = 9'h113 == io_addr ? mem_275 : _GEN_274; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_276 = 9'h114 == io_addr ? mem_276 : _GEN_275; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_277 = 9'h115 == io_addr ? mem_277 : _GEN_276; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_278 = 9'h116 == io_addr ? mem_278 : _GEN_277; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_279 = 9'h117 == io_addr ? mem_279 : _GEN_278; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_280 = 9'h118 == io_addr ? mem_280 : _GEN_279; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_281 = 9'h119 == io_addr ? mem_281 : _GEN_280; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_282 = 9'h11a == io_addr ? mem_282 : _GEN_281; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_283 = 9'h11b == io_addr ? mem_283 : _GEN_282; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_284 = 9'h11c == io_addr ? mem_284 : _GEN_283; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_285 = 9'h11d == io_addr ? mem_285 : _GEN_284; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_286 = 9'h11e == io_addr ? mem_286 : _GEN_285; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_287 = 9'h11f == io_addr ? mem_287 : _GEN_286; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_288 = 9'h120 == io_addr ? mem_288 : _GEN_287; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_289 = 9'h121 == io_addr ? mem_289 : _GEN_288; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_290 = 9'h122 == io_addr ? mem_290 : _GEN_289; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_291 = 9'h123 == io_addr ? mem_291 : _GEN_290; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_292 = 9'h124 == io_addr ? mem_292 : _GEN_291; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_293 = 9'h125 == io_addr ? mem_293 : _GEN_292; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_294 = 9'h126 == io_addr ? mem_294 : _GEN_293; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_295 = 9'h127 == io_addr ? mem_295 : _GEN_294; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_296 = 9'h128 == io_addr ? mem_296 : _GEN_295; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_297 = 9'h129 == io_addr ? mem_297 : _GEN_296; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_298 = 9'h12a == io_addr ? mem_298 : _GEN_297; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_299 = 9'h12b == io_addr ? mem_299 : _GEN_298; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_300 = 9'h12c == io_addr ? mem_300 : _GEN_299; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_301 = 9'h12d == io_addr ? mem_301 : _GEN_300; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_302 = 9'h12e == io_addr ? mem_302 : _GEN_301; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_303 = 9'h12f == io_addr ? mem_303 : _GEN_302; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_304 = 9'h130 == io_addr ? mem_304 : _GEN_303; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_305 = 9'h131 == io_addr ? mem_305 : _GEN_304; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_306 = 9'h132 == io_addr ? mem_306 : _GEN_305; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_307 = 9'h133 == io_addr ? mem_307 : _GEN_306; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_308 = 9'h134 == io_addr ? mem_308 : _GEN_307; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_309 = 9'h135 == io_addr ? mem_309 : _GEN_308; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_310 = 9'h136 == io_addr ? mem_310 : _GEN_309; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_311 = 9'h137 == io_addr ? mem_311 : _GEN_310; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_312 = 9'h138 == io_addr ? mem_312 : _GEN_311; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_313 = 9'h139 == io_addr ? mem_313 : _GEN_312; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_314 = 9'h13a == io_addr ? mem_314 : _GEN_313; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_315 = 9'h13b == io_addr ? mem_315 : _GEN_314; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_316 = 9'h13c == io_addr ? mem_316 : _GEN_315; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_317 = 9'h13d == io_addr ? mem_317 : _GEN_316; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_318 = 9'h13e == io_addr ? mem_318 : _GEN_317; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_319 = 9'h13f == io_addr ? mem_319 : _GEN_318; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_320 = 9'h140 == io_addr ? mem_320 : _GEN_319; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_321 = 9'h141 == io_addr ? mem_321 : _GEN_320; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_322 = 9'h142 == io_addr ? mem_322 : _GEN_321; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_323 = 9'h143 == io_addr ? mem_323 : _GEN_322; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_324 = 9'h144 == io_addr ? mem_324 : _GEN_323; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_325 = 9'h145 == io_addr ? mem_325 : _GEN_324; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_326 = 9'h146 == io_addr ? mem_326 : _GEN_325; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_327 = 9'h147 == io_addr ? mem_327 : _GEN_326; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_328 = 9'h148 == io_addr ? mem_328 : _GEN_327; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_329 = 9'h149 == io_addr ? mem_329 : _GEN_328; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_330 = 9'h14a == io_addr ? mem_330 : _GEN_329; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_331 = 9'h14b == io_addr ? mem_331 : _GEN_330; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_332 = 9'h14c == io_addr ? mem_332 : _GEN_331; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_333 = 9'h14d == io_addr ? mem_333 : _GEN_332; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_334 = 9'h14e == io_addr ? mem_334 : _GEN_333; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_335 = 9'h14f == io_addr ? mem_335 : _GEN_334; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_336 = 9'h150 == io_addr ? mem_336 : _GEN_335; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_337 = 9'h151 == io_addr ? mem_337 : _GEN_336; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_338 = 9'h152 == io_addr ? mem_338 : _GEN_337; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_339 = 9'h153 == io_addr ? mem_339 : _GEN_338; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_340 = 9'h154 == io_addr ? mem_340 : _GEN_339; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_341 = 9'h155 == io_addr ? mem_341 : _GEN_340; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_342 = 9'h156 == io_addr ? mem_342 : _GEN_341; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_343 = 9'h157 == io_addr ? mem_343 : _GEN_342; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_344 = 9'h158 == io_addr ? mem_344 : _GEN_343; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_345 = 9'h159 == io_addr ? mem_345 : _GEN_344; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_346 = 9'h15a == io_addr ? mem_346 : _GEN_345; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_347 = 9'h15b == io_addr ? mem_347 : _GEN_346; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_348 = 9'h15c == io_addr ? mem_348 : _GEN_347; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_349 = 9'h15d == io_addr ? mem_349 : _GEN_348; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_350 = 9'h15e == io_addr ? mem_350 : _GEN_349; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_351 = 9'h15f == io_addr ? mem_351 : _GEN_350; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_352 = 9'h160 == io_addr ? mem_352 : _GEN_351; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_353 = 9'h161 == io_addr ? mem_353 : _GEN_352; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_354 = 9'h162 == io_addr ? mem_354 : _GEN_353; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_355 = 9'h163 == io_addr ? mem_355 : _GEN_354; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_356 = 9'h164 == io_addr ? mem_356 : _GEN_355; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_357 = 9'h165 == io_addr ? mem_357 : _GEN_356; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_358 = 9'h166 == io_addr ? mem_358 : _GEN_357; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_359 = 9'h167 == io_addr ? mem_359 : _GEN_358; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_360 = 9'h168 == io_addr ? mem_360 : _GEN_359; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_361 = 9'h169 == io_addr ? mem_361 : _GEN_360; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_362 = 9'h16a == io_addr ? mem_362 : _GEN_361; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_363 = 9'h16b == io_addr ? mem_363 : _GEN_362; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_364 = 9'h16c == io_addr ? mem_364 : _GEN_363; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_365 = 9'h16d == io_addr ? mem_365 : _GEN_364; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_366 = 9'h16e == io_addr ? mem_366 : _GEN_365; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_367 = 9'h16f == io_addr ? mem_367 : _GEN_366; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_368 = 9'h170 == io_addr ? mem_368 : _GEN_367; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_369 = 9'h171 == io_addr ? mem_369 : _GEN_368; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_370 = 9'h172 == io_addr ? mem_370 : _GEN_369; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_371 = 9'h173 == io_addr ? mem_371 : _GEN_370; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_372 = 9'h174 == io_addr ? mem_372 : _GEN_371; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_373 = 9'h175 == io_addr ? mem_373 : _GEN_372; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_374 = 9'h176 == io_addr ? mem_374 : _GEN_373; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_375 = 9'h177 == io_addr ? mem_375 : _GEN_374; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_376 = 9'h178 == io_addr ? mem_376 : _GEN_375; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_377 = 9'h179 == io_addr ? mem_377 : _GEN_376; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_378 = 9'h17a == io_addr ? mem_378 : _GEN_377; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_379 = 9'h17b == io_addr ? mem_379 : _GEN_378; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_380 = 9'h17c == io_addr ? mem_380 : _GEN_379; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_381 = 9'h17d == io_addr ? mem_381 : _GEN_380; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_382 = 9'h17e == io_addr ? mem_382 : _GEN_381; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_383 = 9'h17f == io_addr ? mem_383 : _GEN_382; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_384 = 9'h180 == io_addr ? mem_384 : _GEN_383; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_385 = 9'h181 == io_addr ? mem_385 : _GEN_384; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_386 = 9'h182 == io_addr ? mem_386 : _GEN_385; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_387 = 9'h183 == io_addr ? mem_387 : _GEN_386; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_388 = 9'h184 == io_addr ? mem_388 : _GEN_387; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_389 = 9'h185 == io_addr ? mem_389 : _GEN_388; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_390 = 9'h186 == io_addr ? mem_390 : _GEN_389; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_391 = 9'h187 == io_addr ? mem_391 : _GEN_390; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_392 = 9'h188 == io_addr ? mem_392 : _GEN_391; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_393 = 9'h189 == io_addr ? mem_393 : _GEN_392; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_394 = 9'h18a == io_addr ? mem_394 : _GEN_393; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_395 = 9'h18b == io_addr ? mem_395 : _GEN_394; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_396 = 9'h18c == io_addr ? mem_396 : _GEN_395; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_397 = 9'h18d == io_addr ? mem_397 : _GEN_396; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_398 = 9'h18e == io_addr ? mem_398 : _GEN_397; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_399 = 9'h18f == io_addr ? mem_399 : _GEN_398; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_400 = 9'h190 == io_addr ? mem_400 : _GEN_399; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_401 = 9'h191 == io_addr ? mem_401 : _GEN_400; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_402 = 9'h192 == io_addr ? mem_402 : _GEN_401; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_403 = 9'h193 == io_addr ? mem_403 : _GEN_402; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_404 = 9'h194 == io_addr ? mem_404 : _GEN_403; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_405 = 9'h195 == io_addr ? mem_405 : _GEN_404; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_406 = 9'h196 == io_addr ? mem_406 : _GEN_405; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_407 = 9'h197 == io_addr ? mem_407 : _GEN_406; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_408 = 9'h198 == io_addr ? mem_408 : _GEN_407; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_409 = 9'h199 == io_addr ? mem_409 : _GEN_408; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_410 = 9'h19a == io_addr ? mem_410 : _GEN_409; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_411 = 9'h19b == io_addr ? mem_411 : _GEN_410; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_412 = 9'h19c == io_addr ? mem_412 : _GEN_411; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_413 = 9'h19d == io_addr ? mem_413 : _GEN_412; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_414 = 9'h19e == io_addr ? mem_414 : _GEN_413; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_415 = 9'h19f == io_addr ? mem_415 : _GEN_414; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_416 = 9'h1a0 == io_addr ? mem_416 : _GEN_415; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_417 = 9'h1a1 == io_addr ? mem_417 : _GEN_416; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_418 = 9'h1a2 == io_addr ? mem_418 : _GEN_417; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_419 = 9'h1a3 == io_addr ? mem_419 : _GEN_418; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_420 = 9'h1a4 == io_addr ? mem_420 : _GEN_419; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_421 = 9'h1a5 == io_addr ? mem_421 : _GEN_420; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_422 = 9'h1a6 == io_addr ? mem_422 : _GEN_421; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_423 = 9'h1a7 == io_addr ? mem_423 : _GEN_422; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_424 = 9'h1a8 == io_addr ? mem_424 : _GEN_423; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_425 = 9'h1a9 == io_addr ? mem_425 : _GEN_424; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_426 = 9'h1aa == io_addr ? mem_426 : _GEN_425; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_427 = 9'h1ab == io_addr ? mem_427 : _GEN_426; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_428 = 9'h1ac == io_addr ? mem_428 : _GEN_427; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_429 = 9'h1ad == io_addr ? mem_429 : _GEN_428; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_430 = 9'h1ae == io_addr ? mem_430 : _GEN_429; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_431 = 9'h1af == io_addr ? mem_431 : _GEN_430; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_432 = 9'h1b0 == io_addr ? mem_432 : _GEN_431; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_433 = 9'h1b1 == io_addr ? mem_433 : _GEN_432; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_434 = 9'h1b2 == io_addr ? mem_434 : _GEN_433; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_435 = 9'h1b3 == io_addr ? mem_435 : _GEN_434; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_436 = 9'h1b4 == io_addr ? mem_436 : _GEN_435; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_437 = 9'h1b5 == io_addr ? mem_437 : _GEN_436; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_438 = 9'h1b6 == io_addr ? mem_438 : _GEN_437; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_439 = 9'h1b7 == io_addr ? mem_439 : _GEN_438; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_440 = 9'h1b8 == io_addr ? mem_440 : _GEN_439; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_441 = 9'h1b9 == io_addr ? mem_441 : _GEN_440; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_442 = 9'h1ba == io_addr ? mem_442 : _GEN_441; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_443 = 9'h1bb == io_addr ? mem_443 : _GEN_442; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_444 = 9'h1bc == io_addr ? mem_444 : _GEN_443; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_445 = 9'h1bd == io_addr ? mem_445 : _GEN_444; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_446 = 9'h1be == io_addr ? mem_446 : _GEN_445; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_447 = 9'h1bf == io_addr ? mem_447 : _GEN_446; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_448 = 9'h1c0 == io_addr ? mem_448 : _GEN_447; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_449 = 9'h1c1 == io_addr ? mem_449 : _GEN_448; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_450 = 9'h1c2 == io_addr ? mem_450 : _GEN_449; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_451 = 9'h1c3 == io_addr ? mem_451 : _GEN_450; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_452 = 9'h1c4 == io_addr ? mem_452 : _GEN_451; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_453 = 9'h1c5 == io_addr ? mem_453 : _GEN_452; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_454 = 9'h1c6 == io_addr ? mem_454 : _GEN_453; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_455 = 9'h1c7 == io_addr ? mem_455 : _GEN_454; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_456 = 9'h1c8 == io_addr ? mem_456 : _GEN_455; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_457 = 9'h1c9 == io_addr ? mem_457 : _GEN_456; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_458 = 9'h1ca == io_addr ? mem_458 : _GEN_457; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_459 = 9'h1cb == io_addr ? mem_459 : _GEN_458; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_460 = 9'h1cc == io_addr ? mem_460 : _GEN_459; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_461 = 9'h1cd == io_addr ? mem_461 : _GEN_460; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_462 = 9'h1ce == io_addr ? mem_462 : _GEN_461; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_463 = 9'h1cf == io_addr ? mem_463 : _GEN_462; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_464 = 9'h1d0 == io_addr ? mem_464 : _GEN_463; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_465 = 9'h1d1 == io_addr ? mem_465 : _GEN_464; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_466 = 9'h1d2 == io_addr ? mem_466 : _GEN_465; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_467 = 9'h1d3 == io_addr ? mem_467 : _GEN_466; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_468 = 9'h1d4 == io_addr ? mem_468 : _GEN_467; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_469 = 9'h1d5 == io_addr ? mem_469 : _GEN_468; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_470 = 9'h1d6 == io_addr ? mem_470 : _GEN_469; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_471 = 9'h1d7 == io_addr ? mem_471 : _GEN_470; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_472 = 9'h1d8 == io_addr ? mem_472 : _GEN_471; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_473 = 9'h1d9 == io_addr ? mem_473 : _GEN_472; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_474 = 9'h1da == io_addr ? mem_474 : _GEN_473; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_475 = 9'h1db == io_addr ? mem_475 : _GEN_474; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_476 = 9'h1dc == io_addr ? mem_476 : _GEN_475; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_477 = 9'h1dd == io_addr ? mem_477 : _GEN_476; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_478 = 9'h1de == io_addr ? mem_478 : _GEN_477; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_479 = 9'h1df == io_addr ? mem_479 : _GEN_478; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_480 = 9'h1e0 == io_addr ? mem_480 : _GEN_479; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_481 = 9'h1e1 == io_addr ? mem_481 : _GEN_480; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_482 = 9'h1e2 == io_addr ? mem_482 : _GEN_481; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_483 = 9'h1e3 == io_addr ? mem_483 : _GEN_482; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_484 = 9'h1e4 == io_addr ? mem_484 : _GEN_483; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_485 = 9'h1e5 == io_addr ? mem_485 : _GEN_484; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_486 = 9'h1e6 == io_addr ? mem_486 : _GEN_485; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_487 = 9'h1e7 == io_addr ? mem_487 : _GEN_486; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_488 = 9'h1e8 == io_addr ? mem_488 : _GEN_487; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_489 = 9'h1e9 == io_addr ? mem_489 : _GEN_488; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_490 = 9'h1ea == io_addr ? mem_490 : _GEN_489; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_491 = 9'h1eb == io_addr ? mem_491 : _GEN_490; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_492 = 9'h1ec == io_addr ? mem_492 : _GEN_491; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_493 = 9'h1ed == io_addr ? mem_493 : _GEN_492; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_494 = 9'h1ee == io_addr ? mem_494 : _GEN_493; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_495 = 9'h1ef == io_addr ? mem_495 : _GEN_494; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_496 = 9'h1f0 == io_addr ? mem_496 : _GEN_495; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_497 = 9'h1f1 == io_addr ? mem_497 : _GEN_496; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_498 = 9'h1f2 == io_addr ? mem_498 : _GEN_497; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_499 = 9'h1f3 == io_addr ? mem_499 : _GEN_498; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_500 = 9'h1f4 == io_addr ? mem_500 : _GEN_499; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_501 = 9'h1f5 == io_addr ? mem_501 : _GEN_500; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_502 = 9'h1f6 == io_addr ? mem_502 : _GEN_501; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_503 = 9'h1f7 == io_addr ? mem_503 : _GEN_502; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_504 = 9'h1f8 == io_addr ? mem_504 : _GEN_503; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_505 = 9'h1f9 == io_addr ? mem_505 : _GEN_504; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_506 = 9'h1fa == io_addr ? mem_506 : _GEN_505; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  wire [18:0] _GEN_507 = 9'h1fb == io_addr ? mem_507 : _GEN_506; // @[RAMWrapper.scala 288:21 RAMWrapper.scala 288:21]
  assign io_dout = io_dout_REG; // @[RAMWrapper.scala 288:11]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_0 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_0 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_1 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_1 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_2 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_2 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_3 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_3 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_4 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_4 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_5 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_5 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_6 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_6 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_7 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_7 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_8 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_8 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_9 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_9 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_10 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_10 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_11 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_11 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_12 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_12 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_13 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_13 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_14 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_14 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_15 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_15 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_16 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_16 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_17 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_17 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_18 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_18 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_19 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_19 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_20 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_20 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_21 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_21 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_22 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_22 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_23 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_23 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_24 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_24 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_25 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_25 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_26 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_26 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_27 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_27 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_28 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_28 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_29 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_29 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_30 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_30 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_31 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_31 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_32 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h20 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_32 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_33 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h21 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_33 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_34 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h22 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_34 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_35 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h23 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_35 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_36 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h24 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_36 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_37 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h25 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_37 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_38 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h26 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_38 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_39 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h27 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_39 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_40 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h28 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_40 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_41 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h29 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_41 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_42 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_42 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_43 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_43 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_44 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_44 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_45 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_45 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_46 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_46 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_47 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h2f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_47 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_48 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h30 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_48 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_49 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h31 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_49 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_50 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h32 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_50 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_51 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h33 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_51 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_52 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h34 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_52 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_53 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h35 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_53 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_54 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h36 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_54 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_55 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h37 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_55 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_56 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h38 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_56 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_57 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h39 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_57 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_58 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_58 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_59 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_59 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_60 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_60 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_61 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_61 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_62 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_62 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_63 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h3f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_63 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_64 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h40 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_64 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_65 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h41 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_65 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_66 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h42 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_66 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_67 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h43 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_67 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_68 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h44 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_68 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_69 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h45 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_69 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_70 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h46 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_70 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_71 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h47 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_71 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_72 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h48 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_72 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_73 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h49 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_73 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_74 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_74 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_75 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_75 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_76 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_76 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_77 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_77 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_78 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_78 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_79 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h4f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_79 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_80 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h50 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_80 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_81 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h51 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_81 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_82 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h52 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_82 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_83 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h53 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_83 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_84 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h54 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_84 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_85 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h55 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_85 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_86 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h56 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_86 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_87 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h57 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_87 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_88 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h58 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_88 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_89 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h59 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_89 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_90 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_90 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_91 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_91 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_92 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_92 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_93 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_93 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_94 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_94 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_95 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h5f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_95 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_96 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h60 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_96 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_97 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h61 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_97 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_98 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h62 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_98 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_99 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h63 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_99 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_100 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h64 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_100 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_101 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h65 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_101 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_102 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h66 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_102 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_103 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h67 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_103 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_104 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h68 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_104 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_105 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h69 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_105 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_106 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_106 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_107 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_107 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_108 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_108 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_109 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_109 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_110 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_110 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_111 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h6f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_111 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_112 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h70 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_112 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_113 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h71 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_113 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_114 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h72 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_114 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_115 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h73 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_115 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_116 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h74 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_116 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_117 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h75 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_117 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_118 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h76 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_118 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_119 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h77 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_119 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_120 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h78 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_120 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_121 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h79 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_121 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_122 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_122 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_123 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_123 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_124 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_124 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_125 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_125 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_126 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_126 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_127 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h7f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_127 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_128 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h80 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_128 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_129 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h81 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_129 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_130 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h82 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_130 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_131 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h83 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_131 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_132 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h84 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_132 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_133 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h85 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_133 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_134 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h86 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_134 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_135 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h87 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_135 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_136 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h88 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_136 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_137 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h89 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_137 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_138 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_138 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_139 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_139 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_140 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_140 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_141 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_141 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_142 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_142 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_143 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h8f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_143 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_144 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h90 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_144 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_145 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h91 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_145 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_146 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h92 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_146 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_147 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h93 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_147 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_148 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h94 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_148 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_149 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h95 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_149 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_150 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h96 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_150 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_151 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h97 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_151 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_152 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h98 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_152 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_153 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h99 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_153 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_154 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_154 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_155 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_155 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_156 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_156 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_157 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_157 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_158 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_158 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_159 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h9f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_159 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_160 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_160 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_161 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_161 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_162 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_162 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_163 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_163 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_164 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_164 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_165 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_165 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_166 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_166 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_167 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_167 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_168 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_168 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_169 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'ha9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_169 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_170 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'haa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_170 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_171 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hab == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_171 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_172 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hac == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_172 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_173 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'had == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_173 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_174 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hae == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_174 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_175 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'haf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_175 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_176 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_176 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_177 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_177 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_178 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_178 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_179 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_179 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_180 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_180 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_181 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_181 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_182 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_182 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_183 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_183 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_184 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_184 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_185 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hb9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_185 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_186 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hba == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_186 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_187 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_187 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_188 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_188 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_189 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_189 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_190 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_190 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_191 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hbf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_191 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_192 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_192 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_193 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_193 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_194 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_194 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_195 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_195 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_196 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_196 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_197 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_197 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_198 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_198 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_199 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_199 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_200 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_200 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_201 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hc9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_201 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_202 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hca == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_202 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_203 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_203 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_204 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_204 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_205 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_205 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_206 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hce == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_206 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_207 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hcf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_207 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_208 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_208 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_209 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_209 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_210 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_210 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_211 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_211 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_212 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_212 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_213 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_213 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_214 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_214 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_215 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_215 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_216 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_216 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_217 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hd9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_217 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_218 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hda == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_218 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_219 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_219 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_220 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_220 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_221 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_221 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_222 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hde == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_222 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_223 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hdf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_223 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_224 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_224 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_225 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_225 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_226 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_226 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_227 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_227 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_228 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_228 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_229 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_229 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_230 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_230 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_231 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_231 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_232 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_232 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_233 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'he9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_233 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_234 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hea == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_234 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_235 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'heb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_235 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_236 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hec == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_236 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_237 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hed == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_237 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_238 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hee == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_238 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_239 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hef == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_239 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_240 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_240 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_241 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_241 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_242 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_242 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_243 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_243 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_244 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_244 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_245 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_245 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_246 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_246 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_247 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_247 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_248 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_248 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_249 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hf9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_249 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_250 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_250 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_251 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_251 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_252 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_252 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_253 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_253 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_254 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hfe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_254 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_255 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'hff == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_255 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_256 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h100 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_256 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_257 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h101 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_257 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_258 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h102 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_258 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_259 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h103 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_259 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_260 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h104 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_260 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_261 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h105 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_261 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_262 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h106 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_262 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_263 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h107 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_263 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_264 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h108 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_264 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_265 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h109 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_265 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_266 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_266 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_267 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_267 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_268 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_268 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_269 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_269 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_270 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_270 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_271 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h10f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_271 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_272 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h110 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_272 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_273 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h111 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_273 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_274 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h112 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_274 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_275 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h113 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_275 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_276 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h114 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_276 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_277 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h115 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_277 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_278 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h116 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_278 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_279 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h117 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_279 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_280 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h118 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_280 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_281 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h119 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_281 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_282 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_282 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_283 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_283 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_284 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_284 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_285 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_285 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_286 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_286 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_287 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h11f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_287 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_288 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h120 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_288 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_289 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h121 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_289 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_290 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h122 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_290 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_291 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h123 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_291 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_292 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h124 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_292 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_293 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h125 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_293 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_294 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h126 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_294 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_295 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h127 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_295 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_296 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h128 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_296 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_297 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h129 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_297 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_298 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_298 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_299 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_299 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_300 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_300 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_301 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_301 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_302 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_302 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_303 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h12f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_303 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_304 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h130 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_304 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_305 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h131 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_305 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_306 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h132 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_306 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_307 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h133 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_307 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_308 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h134 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_308 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_309 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h135 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_309 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_310 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h136 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_310 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_311 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h137 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_311 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_312 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h138 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_312 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_313 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h139 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_313 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_314 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_314 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_315 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_315 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_316 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_316 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_317 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_317 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_318 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_318 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_319 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h13f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_319 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_320 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h140 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_320 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_321 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h141 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_321 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_322 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h142 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_322 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_323 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h143 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_323 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_324 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h144 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_324 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_325 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h145 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_325 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_326 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h146 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_326 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_327 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h147 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_327 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_328 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h148 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_328 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_329 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h149 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_329 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_330 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_330 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_331 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_331 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_332 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_332 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_333 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_333 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_334 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_334 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_335 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h14f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_335 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_336 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h150 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_336 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_337 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h151 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_337 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_338 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h152 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_338 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_339 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h153 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_339 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_340 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h154 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_340 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_341 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h155 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_341 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_342 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h156 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_342 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_343 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h157 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_343 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_344 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h158 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_344 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_345 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h159 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_345 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_346 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_346 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_347 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_347 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_348 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_348 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_349 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_349 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_350 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_350 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_351 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h15f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_351 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_352 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h160 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_352 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_353 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h161 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_353 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_354 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h162 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_354 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_355 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h163 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_355 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_356 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h164 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_356 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_357 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h165 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_357 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_358 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h166 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_358 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_359 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h167 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_359 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_360 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h168 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_360 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_361 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h169 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_361 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_362 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_362 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_363 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_363 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_364 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_364 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_365 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_365 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_366 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_366 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_367 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h16f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_367 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_368 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h170 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_368 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_369 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h171 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_369 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_370 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h172 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_370 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_371 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h173 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_371 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_372 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h174 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_372 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_373 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h175 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_373 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_374 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h176 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_374 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_375 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h177 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_375 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_376 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h178 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_376 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_377 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h179 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_377 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_378 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_378 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_379 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_379 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_380 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_380 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_381 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_381 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_382 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_382 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_383 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h17f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_383 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_384 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h180 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_384 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_385 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h181 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_385 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_386 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h182 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_386 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_387 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h183 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_387 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_388 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h184 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_388 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_389 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h185 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_389 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_390 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h186 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_390 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_391 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h187 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_391 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_392 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h188 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_392 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_393 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h189 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_393 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_394 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_394 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_395 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_395 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_396 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_396 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_397 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_397 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_398 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_398 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_399 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h18f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_399 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_400 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h190 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_400 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_401 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h191 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_401 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_402 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h192 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_402 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_403 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h193 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_403 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_404 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h194 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_404 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_405 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h195 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_405 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_406 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h196 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_406 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_407 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h197 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_407 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_408 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h198 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_408 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_409 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h199 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_409 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_410 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19a == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_410 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_411 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19b == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_411 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_412 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19c == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_412 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_413 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19d == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_413 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_414 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19e == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_414 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_415 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h19f == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_415 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_416 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_416 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_417 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_417 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_418 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_418 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_419 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_419 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_420 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_420 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_421 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_421 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_422 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_422 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_423 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_423 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_424 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_424 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_425 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1a9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_425 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_426 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1aa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_426 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_427 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ab == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_427 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_428 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ac == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_428 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_429 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ad == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_429 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_430 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ae == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_430 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_431 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1af == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_431 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_432 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_432 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_433 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_433 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_434 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_434 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_435 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_435 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_436 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_436 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_437 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_437 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_438 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_438 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_439 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_439 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_440 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_440 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_441 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1b9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_441 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_442 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ba == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_442 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_443 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_443 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_444 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_444 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_445 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_445 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_446 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1be == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_446 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_447 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1bf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_447 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_448 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_448 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_449 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_449 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_450 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_450 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_451 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_451 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_452 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_452 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_453 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_453 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_454 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_454 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_455 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_455 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_456 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_456 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_457 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1c9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_457 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_458 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ca == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_458 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_459 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_459 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_460 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_460 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_461 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_461 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_462 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ce == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_462 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_463 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1cf == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_463 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_464 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_464 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_465 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_465 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_466 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_466 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_467 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_467 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_468 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_468 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_469 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_469 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_470 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_470 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_471 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_471 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_472 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_472 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_473 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1d9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_473 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_474 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1da == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_474 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_475 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1db == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_475 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_476 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1dc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_476 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_477 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1dd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_477 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_478 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1de == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_478 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_479 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1df == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_479 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_480 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_480 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_481 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_481 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_482 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_482 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_483 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_483 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_484 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_484 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_485 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_485 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_486 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_486 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_487 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_487 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_488 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_488 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_489 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1e9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_489 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_490 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ea == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_490 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_491 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1eb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_491 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_492 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ec == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_492 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_493 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ed == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_493 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_494 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ee == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_494 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_495 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ef == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_495 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_496 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f0 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_496 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_497 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f1 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_497 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_498 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f2 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_498 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_499 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f3 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_499 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_500 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f4 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_500 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_501 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f5 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_501 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_502 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f6 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_502 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_503 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f7 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_503 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_504 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f8 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_504 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_505 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1f9 == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_505 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_506 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fa == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_506 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_507 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fb == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_507 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_508 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fc == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_508 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_509 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fd == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_509 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_510 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1fe == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_510 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 286:20]
      mem_511 <= 19'h0; // @[RAMWrapper.scala 286:20]
    end else if (io_we) begin // @[RAMWrapper.scala 290:15]
      if (9'h1ff == io_addr) begin // @[RAMWrapper.scala 291:18]
        mem_511 <= io_din; // @[RAMWrapper.scala 291:18]
      end
    end
    if (9'h1ff == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_511; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fe == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_510; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fd == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_509; // @[RAMWrapper.scala 288:21]
    end else if (9'h1fc == io_addr) begin // @[RAMWrapper.scala 288:21]
      io_dout_REG <= mem_508; // @[RAMWrapper.scala 288:21]
    end else begin
      io_dout_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[18:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[18:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[18:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[18:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[18:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[18:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[18:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[18:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[18:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[18:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[18:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[18:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[18:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[18:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[18:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[18:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[18:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[18:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[18:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[18:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[18:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[18:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[18:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[18:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[18:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[18:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[18:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[18:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[18:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[18:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[18:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[18:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[18:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[18:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[18:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[18:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[18:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[18:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[18:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[18:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[18:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[18:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[18:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[18:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[18:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[18:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[18:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[18:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[18:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[18:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[18:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[18:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[18:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[18:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[18:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[18:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[18:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[18:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[18:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[18:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[18:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[18:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[18:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[18:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[18:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[18:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[18:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[18:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[18:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[18:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[18:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[18:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[18:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[18:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[18:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[18:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[18:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[18:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[18:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[18:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[18:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[18:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[18:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[18:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[18:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[18:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[18:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[18:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[18:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[18:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[18:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[18:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[18:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[18:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[18:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[18:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[18:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[18:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[18:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[18:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[18:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[18:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[18:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[18:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[18:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[18:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[18:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[18:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[18:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[18:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[18:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[18:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[18:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[18:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[18:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[18:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[18:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[18:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[18:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[18:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[18:0];
  _RAND_128 = {1{`RANDOM}};
  mem_128 = _RAND_128[18:0];
  _RAND_129 = {1{`RANDOM}};
  mem_129 = _RAND_129[18:0];
  _RAND_130 = {1{`RANDOM}};
  mem_130 = _RAND_130[18:0];
  _RAND_131 = {1{`RANDOM}};
  mem_131 = _RAND_131[18:0];
  _RAND_132 = {1{`RANDOM}};
  mem_132 = _RAND_132[18:0];
  _RAND_133 = {1{`RANDOM}};
  mem_133 = _RAND_133[18:0];
  _RAND_134 = {1{`RANDOM}};
  mem_134 = _RAND_134[18:0];
  _RAND_135 = {1{`RANDOM}};
  mem_135 = _RAND_135[18:0];
  _RAND_136 = {1{`RANDOM}};
  mem_136 = _RAND_136[18:0];
  _RAND_137 = {1{`RANDOM}};
  mem_137 = _RAND_137[18:0];
  _RAND_138 = {1{`RANDOM}};
  mem_138 = _RAND_138[18:0];
  _RAND_139 = {1{`RANDOM}};
  mem_139 = _RAND_139[18:0];
  _RAND_140 = {1{`RANDOM}};
  mem_140 = _RAND_140[18:0];
  _RAND_141 = {1{`RANDOM}};
  mem_141 = _RAND_141[18:0];
  _RAND_142 = {1{`RANDOM}};
  mem_142 = _RAND_142[18:0];
  _RAND_143 = {1{`RANDOM}};
  mem_143 = _RAND_143[18:0];
  _RAND_144 = {1{`RANDOM}};
  mem_144 = _RAND_144[18:0];
  _RAND_145 = {1{`RANDOM}};
  mem_145 = _RAND_145[18:0];
  _RAND_146 = {1{`RANDOM}};
  mem_146 = _RAND_146[18:0];
  _RAND_147 = {1{`RANDOM}};
  mem_147 = _RAND_147[18:0];
  _RAND_148 = {1{`RANDOM}};
  mem_148 = _RAND_148[18:0];
  _RAND_149 = {1{`RANDOM}};
  mem_149 = _RAND_149[18:0];
  _RAND_150 = {1{`RANDOM}};
  mem_150 = _RAND_150[18:0];
  _RAND_151 = {1{`RANDOM}};
  mem_151 = _RAND_151[18:0];
  _RAND_152 = {1{`RANDOM}};
  mem_152 = _RAND_152[18:0];
  _RAND_153 = {1{`RANDOM}};
  mem_153 = _RAND_153[18:0];
  _RAND_154 = {1{`RANDOM}};
  mem_154 = _RAND_154[18:0];
  _RAND_155 = {1{`RANDOM}};
  mem_155 = _RAND_155[18:0];
  _RAND_156 = {1{`RANDOM}};
  mem_156 = _RAND_156[18:0];
  _RAND_157 = {1{`RANDOM}};
  mem_157 = _RAND_157[18:0];
  _RAND_158 = {1{`RANDOM}};
  mem_158 = _RAND_158[18:0];
  _RAND_159 = {1{`RANDOM}};
  mem_159 = _RAND_159[18:0];
  _RAND_160 = {1{`RANDOM}};
  mem_160 = _RAND_160[18:0];
  _RAND_161 = {1{`RANDOM}};
  mem_161 = _RAND_161[18:0];
  _RAND_162 = {1{`RANDOM}};
  mem_162 = _RAND_162[18:0];
  _RAND_163 = {1{`RANDOM}};
  mem_163 = _RAND_163[18:0];
  _RAND_164 = {1{`RANDOM}};
  mem_164 = _RAND_164[18:0];
  _RAND_165 = {1{`RANDOM}};
  mem_165 = _RAND_165[18:0];
  _RAND_166 = {1{`RANDOM}};
  mem_166 = _RAND_166[18:0];
  _RAND_167 = {1{`RANDOM}};
  mem_167 = _RAND_167[18:0];
  _RAND_168 = {1{`RANDOM}};
  mem_168 = _RAND_168[18:0];
  _RAND_169 = {1{`RANDOM}};
  mem_169 = _RAND_169[18:0];
  _RAND_170 = {1{`RANDOM}};
  mem_170 = _RAND_170[18:0];
  _RAND_171 = {1{`RANDOM}};
  mem_171 = _RAND_171[18:0];
  _RAND_172 = {1{`RANDOM}};
  mem_172 = _RAND_172[18:0];
  _RAND_173 = {1{`RANDOM}};
  mem_173 = _RAND_173[18:0];
  _RAND_174 = {1{`RANDOM}};
  mem_174 = _RAND_174[18:0];
  _RAND_175 = {1{`RANDOM}};
  mem_175 = _RAND_175[18:0];
  _RAND_176 = {1{`RANDOM}};
  mem_176 = _RAND_176[18:0];
  _RAND_177 = {1{`RANDOM}};
  mem_177 = _RAND_177[18:0];
  _RAND_178 = {1{`RANDOM}};
  mem_178 = _RAND_178[18:0];
  _RAND_179 = {1{`RANDOM}};
  mem_179 = _RAND_179[18:0];
  _RAND_180 = {1{`RANDOM}};
  mem_180 = _RAND_180[18:0];
  _RAND_181 = {1{`RANDOM}};
  mem_181 = _RAND_181[18:0];
  _RAND_182 = {1{`RANDOM}};
  mem_182 = _RAND_182[18:0];
  _RAND_183 = {1{`RANDOM}};
  mem_183 = _RAND_183[18:0];
  _RAND_184 = {1{`RANDOM}};
  mem_184 = _RAND_184[18:0];
  _RAND_185 = {1{`RANDOM}};
  mem_185 = _RAND_185[18:0];
  _RAND_186 = {1{`RANDOM}};
  mem_186 = _RAND_186[18:0];
  _RAND_187 = {1{`RANDOM}};
  mem_187 = _RAND_187[18:0];
  _RAND_188 = {1{`RANDOM}};
  mem_188 = _RAND_188[18:0];
  _RAND_189 = {1{`RANDOM}};
  mem_189 = _RAND_189[18:0];
  _RAND_190 = {1{`RANDOM}};
  mem_190 = _RAND_190[18:0];
  _RAND_191 = {1{`RANDOM}};
  mem_191 = _RAND_191[18:0];
  _RAND_192 = {1{`RANDOM}};
  mem_192 = _RAND_192[18:0];
  _RAND_193 = {1{`RANDOM}};
  mem_193 = _RAND_193[18:0];
  _RAND_194 = {1{`RANDOM}};
  mem_194 = _RAND_194[18:0];
  _RAND_195 = {1{`RANDOM}};
  mem_195 = _RAND_195[18:0];
  _RAND_196 = {1{`RANDOM}};
  mem_196 = _RAND_196[18:0];
  _RAND_197 = {1{`RANDOM}};
  mem_197 = _RAND_197[18:0];
  _RAND_198 = {1{`RANDOM}};
  mem_198 = _RAND_198[18:0];
  _RAND_199 = {1{`RANDOM}};
  mem_199 = _RAND_199[18:0];
  _RAND_200 = {1{`RANDOM}};
  mem_200 = _RAND_200[18:0];
  _RAND_201 = {1{`RANDOM}};
  mem_201 = _RAND_201[18:0];
  _RAND_202 = {1{`RANDOM}};
  mem_202 = _RAND_202[18:0];
  _RAND_203 = {1{`RANDOM}};
  mem_203 = _RAND_203[18:0];
  _RAND_204 = {1{`RANDOM}};
  mem_204 = _RAND_204[18:0];
  _RAND_205 = {1{`RANDOM}};
  mem_205 = _RAND_205[18:0];
  _RAND_206 = {1{`RANDOM}};
  mem_206 = _RAND_206[18:0];
  _RAND_207 = {1{`RANDOM}};
  mem_207 = _RAND_207[18:0];
  _RAND_208 = {1{`RANDOM}};
  mem_208 = _RAND_208[18:0];
  _RAND_209 = {1{`RANDOM}};
  mem_209 = _RAND_209[18:0];
  _RAND_210 = {1{`RANDOM}};
  mem_210 = _RAND_210[18:0];
  _RAND_211 = {1{`RANDOM}};
  mem_211 = _RAND_211[18:0];
  _RAND_212 = {1{`RANDOM}};
  mem_212 = _RAND_212[18:0];
  _RAND_213 = {1{`RANDOM}};
  mem_213 = _RAND_213[18:0];
  _RAND_214 = {1{`RANDOM}};
  mem_214 = _RAND_214[18:0];
  _RAND_215 = {1{`RANDOM}};
  mem_215 = _RAND_215[18:0];
  _RAND_216 = {1{`RANDOM}};
  mem_216 = _RAND_216[18:0];
  _RAND_217 = {1{`RANDOM}};
  mem_217 = _RAND_217[18:0];
  _RAND_218 = {1{`RANDOM}};
  mem_218 = _RAND_218[18:0];
  _RAND_219 = {1{`RANDOM}};
  mem_219 = _RAND_219[18:0];
  _RAND_220 = {1{`RANDOM}};
  mem_220 = _RAND_220[18:0];
  _RAND_221 = {1{`RANDOM}};
  mem_221 = _RAND_221[18:0];
  _RAND_222 = {1{`RANDOM}};
  mem_222 = _RAND_222[18:0];
  _RAND_223 = {1{`RANDOM}};
  mem_223 = _RAND_223[18:0];
  _RAND_224 = {1{`RANDOM}};
  mem_224 = _RAND_224[18:0];
  _RAND_225 = {1{`RANDOM}};
  mem_225 = _RAND_225[18:0];
  _RAND_226 = {1{`RANDOM}};
  mem_226 = _RAND_226[18:0];
  _RAND_227 = {1{`RANDOM}};
  mem_227 = _RAND_227[18:0];
  _RAND_228 = {1{`RANDOM}};
  mem_228 = _RAND_228[18:0];
  _RAND_229 = {1{`RANDOM}};
  mem_229 = _RAND_229[18:0];
  _RAND_230 = {1{`RANDOM}};
  mem_230 = _RAND_230[18:0];
  _RAND_231 = {1{`RANDOM}};
  mem_231 = _RAND_231[18:0];
  _RAND_232 = {1{`RANDOM}};
  mem_232 = _RAND_232[18:0];
  _RAND_233 = {1{`RANDOM}};
  mem_233 = _RAND_233[18:0];
  _RAND_234 = {1{`RANDOM}};
  mem_234 = _RAND_234[18:0];
  _RAND_235 = {1{`RANDOM}};
  mem_235 = _RAND_235[18:0];
  _RAND_236 = {1{`RANDOM}};
  mem_236 = _RAND_236[18:0];
  _RAND_237 = {1{`RANDOM}};
  mem_237 = _RAND_237[18:0];
  _RAND_238 = {1{`RANDOM}};
  mem_238 = _RAND_238[18:0];
  _RAND_239 = {1{`RANDOM}};
  mem_239 = _RAND_239[18:0];
  _RAND_240 = {1{`RANDOM}};
  mem_240 = _RAND_240[18:0];
  _RAND_241 = {1{`RANDOM}};
  mem_241 = _RAND_241[18:0];
  _RAND_242 = {1{`RANDOM}};
  mem_242 = _RAND_242[18:0];
  _RAND_243 = {1{`RANDOM}};
  mem_243 = _RAND_243[18:0];
  _RAND_244 = {1{`RANDOM}};
  mem_244 = _RAND_244[18:0];
  _RAND_245 = {1{`RANDOM}};
  mem_245 = _RAND_245[18:0];
  _RAND_246 = {1{`RANDOM}};
  mem_246 = _RAND_246[18:0];
  _RAND_247 = {1{`RANDOM}};
  mem_247 = _RAND_247[18:0];
  _RAND_248 = {1{`RANDOM}};
  mem_248 = _RAND_248[18:0];
  _RAND_249 = {1{`RANDOM}};
  mem_249 = _RAND_249[18:0];
  _RAND_250 = {1{`RANDOM}};
  mem_250 = _RAND_250[18:0];
  _RAND_251 = {1{`RANDOM}};
  mem_251 = _RAND_251[18:0];
  _RAND_252 = {1{`RANDOM}};
  mem_252 = _RAND_252[18:0];
  _RAND_253 = {1{`RANDOM}};
  mem_253 = _RAND_253[18:0];
  _RAND_254 = {1{`RANDOM}};
  mem_254 = _RAND_254[18:0];
  _RAND_255 = {1{`RANDOM}};
  mem_255 = _RAND_255[18:0];
  _RAND_256 = {1{`RANDOM}};
  mem_256 = _RAND_256[18:0];
  _RAND_257 = {1{`RANDOM}};
  mem_257 = _RAND_257[18:0];
  _RAND_258 = {1{`RANDOM}};
  mem_258 = _RAND_258[18:0];
  _RAND_259 = {1{`RANDOM}};
  mem_259 = _RAND_259[18:0];
  _RAND_260 = {1{`RANDOM}};
  mem_260 = _RAND_260[18:0];
  _RAND_261 = {1{`RANDOM}};
  mem_261 = _RAND_261[18:0];
  _RAND_262 = {1{`RANDOM}};
  mem_262 = _RAND_262[18:0];
  _RAND_263 = {1{`RANDOM}};
  mem_263 = _RAND_263[18:0];
  _RAND_264 = {1{`RANDOM}};
  mem_264 = _RAND_264[18:0];
  _RAND_265 = {1{`RANDOM}};
  mem_265 = _RAND_265[18:0];
  _RAND_266 = {1{`RANDOM}};
  mem_266 = _RAND_266[18:0];
  _RAND_267 = {1{`RANDOM}};
  mem_267 = _RAND_267[18:0];
  _RAND_268 = {1{`RANDOM}};
  mem_268 = _RAND_268[18:0];
  _RAND_269 = {1{`RANDOM}};
  mem_269 = _RAND_269[18:0];
  _RAND_270 = {1{`RANDOM}};
  mem_270 = _RAND_270[18:0];
  _RAND_271 = {1{`RANDOM}};
  mem_271 = _RAND_271[18:0];
  _RAND_272 = {1{`RANDOM}};
  mem_272 = _RAND_272[18:0];
  _RAND_273 = {1{`RANDOM}};
  mem_273 = _RAND_273[18:0];
  _RAND_274 = {1{`RANDOM}};
  mem_274 = _RAND_274[18:0];
  _RAND_275 = {1{`RANDOM}};
  mem_275 = _RAND_275[18:0];
  _RAND_276 = {1{`RANDOM}};
  mem_276 = _RAND_276[18:0];
  _RAND_277 = {1{`RANDOM}};
  mem_277 = _RAND_277[18:0];
  _RAND_278 = {1{`RANDOM}};
  mem_278 = _RAND_278[18:0];
  _RAND_279 = {1{`RANDOM}};
  mem_279 = _RAND_279[18:0];
  _RAND_280 = {1{`RANDOM}};
  mem_280 = _RAND_280[18:0];
  _RAND_281 = {1{`RANDOM}};
  mem_281 = _RAND_281[18:0];
  _RAND_282 = {1{`RANDOM}};
  mem_282 = _RAND_282[18:0];
  _RAND_283 = {1{`RANDOM}};
  mem_283 = _RAND_283[18:0];
  _RAND_284 = {1{`RANDOM}};
  mem_284 = _RAND_284[18:0];
  _RAND_285 = {1{`RANDOM}};
  mem_285 = _RAND_285[18:0];
  _RAND_286 = {1{`RANDOM}};
  mem_286 = _RAND_286[18:0];
  _RAND_287 = {1{`RANDOM}};
  mem_287 = _RAND_287[18:0];
  _RAND_288 = {1{`RANDOM}};
  mem_288 = _RAND_288[18:0];
  _RAND_289 = {1{`RANDOM}};
  mem_289 = _RAND_289[18:0];
  _RAND_290 = {1{`RANDOM}};
  mem_290 = _RAND_290[18:0];
  _RAND_291 = {1{`RANDOM}};
  mem_291 = _RAND_291[18:0];
  _RAND_292 = {1{`RANDOM}};
  mem_292 = _RAND_292[18:0];
  _RAND_293 = {1{`RANDOM}};
  mem_293 = _RAND_293[18:0];
  _RAND_294 = {1{`RANDOM}};
  mem_294 = _RAND_294[18:0];
  _RAND_295 = {1{`RANDOM}};
  mem_295 = _RAND_295[18:0];
  _RAND_296 = {1{`RANDOM}};
  mem_296 = _RAND_296[18:0];
  _RAND_297 = {1{`RANDOM}};
  mem_297 = _RAND_297[18:0];
  _RAND_298 = {1{`RANDOM}};
  mem_298 = _RAND_298[18:0];
  _RAND_299 = {1{`RANDOM}};
  mem_299 = _RAND_299[18:0];
  _RAND_300 = {1{`RANDOM}};
  mem_300 = _RAND_300[18:0];
  _RAND_301 = {1{`RANDOM}};
  mem_301 = _RAND_301[18:0];
  _RAND_302 = {1{`RANDOM}};
  mem_302 = _RAND_302[18:0];
  _RAND_303 = {1{`RANDOM}};
  mem_303 = _RAND_303[18:0];
  _RAND_304 = {1{`RANDOM}};
  mem_304 = _RAND_304[18:0];
  _RAND_305 = {1{`RANDOM}};
  mem_305 = _RAND_305[18:0];
  _RAND_306 = {1{`RANDOM}};
  mem_306 = _RAND_306[18:0];
  _RAND_307 = {1{`RANDOM}};
  mem_307 = _RAND_307[18:0];
  _RAND_308 = {1{`RANDOM}};
  mem_308 = _RAND_308[18:0];
  _RAND_309 = {1{`RANDOM}};
  mem_309 = _RAND_309[18:0];
  _RAND_310 = {1{`RANDOM}};
  mem_310 = _RAND_310[18:0];
  _RAND_311 = {1{`RANDOM}};
  mem_311 = _RAND_311[18:0];
  _RAND_312 = {1{`RANDOM}};
  mem_312 = _RAND_312[18:0];
  _RAND_313 = {1{`RANDOM}};
  mem_313 = _RAND_313[18:0];
  _RAND_314 = {1{`RANDOM}};
  mem_314 = _RAND_314[18:0];
  _RAND_315 = {1{`RANDOM}};
  mem_315 = _RAND_315[18:0];
  _RAND_316 = {1{`RANDOM}};
  mem_316 = _RAND_316[18:0];
  _RAND_317 = {1{`RANDOM}};
  mem_317 = _RAND_317[18:0];
  _RAND_318 = {1{`RANDOM}};
  mem_318 = _RAND_318[18:0];
  _RAND_319 = {1{`RANDOM}};
  mem_319 = _RAND_319[18:0];
  _RAND_320 = {1{`RANDOM}};
  mem_320 = _RAND_320[18:0];
  _RAND_321 = {1{`RANDOM}};
  mem_321 = _RAND_321[18:0];
  _RAND_322 = {1{`RANDOM}};
  mem_322 = _RAND_322[18:0];
  _RAND_323 = {1{`RANDOM}};
  mem_323 = _RAND_323[18:0];
  _RAND_324 = {1{`RANDOM}};
  mem_324 = _RAND_324[18:0];
  _RAND_325 = {1{`RANDOM}};
  mem_325 = _RAND_325[18:0];
  _RAND_326 = {1{`RANDOM}};
  mem_326 = _RAND_326[18:0];
  _RAND_327 = {1{`RANDOM}};
  mem_327 = _RAND_327[18:0];
  _RAND_328 = {1{`RANDOM}};
  mem_328 = _RAND_328[18:0];
  _RAND_329 = {1{`RANDOM}};
  mem_329 = _RAND_329[18:0];
  _RAND_330 = {1{`RANDOM}};
  mem_330 = _RAND_330[18:0];
  _RAND_331 = {1{`RANDOM}};
  mem_331 = _RAND_331[18:0];
  _RAND_332 = {1{`RANDOM}};
  mem_332 = _RAND_332[18:0];
  _RAND_333 = {1{`RANDOM}};
  mem_333 = _RAND_333[18:0];
  _RAND_334 = {1{`RANDOM}};
  mem_334 = _RAND_334[18:0];
  _RAND_335 = {1{`RANDOM}};
  mem_335 = _RAND_335[18:0];
  _RAND_336 = {1{`RANDOM}};
  mem_336 = _RAND_336[18:0];
  _RAND_337 = {1{`RANDOM}};
  mem_337 = _RAND_337[18:0];
  _RAND_338 = {1{`RANDOM}};
  mem_338 = _RAND_338[18:0];
  _RAND_339 = {1{`RANDOM}};
  mem_339 = _RAND_339[18:0];
  _RAND_340 = {1{`RANDOM}};
  mem_340 = _RAND_340[18:0];
  _RAND_341 = {1{`RANDOM}};
  mem_341 = _RAND_341[18:0];
  _RAND_342 = {1{`RANDOM}};
  mem_342 = _RAND_342[18:0];
  _RAND_343 = {1{`RANDOM}};
  mem_343 = _RAND_343[18:0];
  _RAND_344 = {1{`RANDOM}};
  mem_344 = _RAND_344[18:0];
  _RAND_345 = {1{`RANDOM}};
  mem_345 = _RAND_345[18:0];
  _RAND_346 = {1{`RANDOM}};
  mem_346 = _RAND_346[18:0];
  _RAND_347 = {1{`RANDOM}};
  mem_347 = _RAND_347[18:0];
  _RAND_348 = {1{`RANDOM}};
  mem_348 = _RAND_348[18:0];
  _RAND_349 = {1{`RANDOM}};
  mem_349 = _RAND_349[18:0];
  _RAND_350 = {1{`RANDOM}};
  mem_350 = _RAND_350[18:0];
  _RAND_351 = {1{`RANDOM}};
  mem_351 = _RAND_351[18:0];
  _RAND_352 = {1{`RANDOM}};
  mem_352 = _RAND_352[18:0];
  _RAND_353 = {1{`RANDOM}};
  mem_353 = _RAND_353[18:0];
  _RAND_354 = {1{`RANDOM}};
  mem_354 = _RAND_354[18:0];
  _RAND_355 = {1{`RANDOM}};
  mem_355 = _RAND_355[18:0];
  _RAND_356 = {1{`RANDOM}};
  mem_356 = _RAND_356[18:0];
  _RAND_357 = {1{`RANDOM}};
  mem_357 = _RAND_357[18:0];
  _RAND_358 = {1{`RANDOM}};
  mem_358 = _RAND_358[18:0];
  _RAND_359 = {1{`RANDOM}};
  mem_359 = _RAND_359[18:0];
  _RAND_360 = {1{`RANDOM}};
  mem_360 = _RAND_360[18:0];
  _RAND_361 = {1{`RANDOM}};
  mem_361 = _RAND_361[18:0];
  _RAND_362 = {1{`RANDOM}};
  mem_362 = _RAND_362[18:0];
  _RAND_363 = {1{`RANDOM}};
  mem_363 = _RAND_363[18:0];
  _RAND_364 = {1{`RANDOM}};
  mem_364 = _RAND_364[18:0];
  _RAND_365 = {1{`RANDOM}};
  mem_365 = _RAND_365[18:0];
  _RAND_366 = {1{`RANDOM}};
  mem_366 = _RAND_366[18:0];
  _RAND_367 = {1{`RANDOM}};
  mem_367 = _RAND_367[18:0];
  _RAND_368 = {1{`RANDOM}};
  mem_368 = _RAND_368[18:0];
  _RAND_369 = {1{`RANDOM}};
  mem_369 = _RAND_369[18:0];
  _RAND_370 = {1{`RANDOM}};
  mem_370 = _RAND_370[18:0];
  _RAND_371 = {1{`RANDOM}};
  mem_371 = _RAND_371[18:0];
  _RAND_372 = {1{`RANDOM}};
  mem_372 = _RAND_372[18:0];
  _RAND_373 = {1{`RANDOM}};
  mem_373 = _RAND_373[18:0];
  _RAND_374 = {1{`RANDOM}};
  mem_374 = _RAND_374[18:0];
  _RAND_375 = {1{`RANDOM}};
  mem_375 = _RAND_375[18:0];
  _RAND_376 = {1{`RANDOM}};
  mem_376 = _RAND_376[18:0];
  _RAND_377 = {1{`RANDOM}};
  mem_377 = _RAND_377[18:0];
  _RAND_378 = {1{`RANDOM}};
  mem_378 = _RAND_378[18:0];
  _RAND_379 = {1{`RANDOM}};
  mem_379 = _RAND_379[18:0];
  _RAND_380 = {1{`RANDOM}};
  mem_380 = _RAND_380[18:0];
  _RAND_381 = {1{`RANDOM}};
  mem_381 = _RAND_381[18:0];
  _RAND_382 = {1{`RANDOM}};
  mem_382 = _RAND_382[18:0];
  _RAND_383 = {1{`RANDOM}};
  mem_383 = _RAND_383[18:0];
  _RAND_384 = {1{`RANDOM}};
  mem_384 = _RAND_384[18:0];
  _RAND_385 = {1{`RANDOM}};
  mem_385 = _RAND_385[18:0];
  _RAND_386 = {1{`RANDOM}};
  mem_386 = _RAND_386[18:0];
  _RAND_387 = {1{`RANDOM}};
  mem_387 = _RAND_387[18:0];
  _RAND_388 = {1{`RANDOM}};
  mem_388 = _RAND_388[18:0];
  _RAND_389 = {1{`RANDOM}};
  mem_389 = _RAND_389[18:0];
  _RAND_390 = {1{`RANDOM}};
  mem_390 = _RAND_390[18:0];
  _RAND_391 = {1{`RANDOM}};
  mem_391 = _RAND_391[18:0];
  _RAND_392 = {1{`RANDOM}};
  mem_392 = _RAND_392[18:0];
  _RAND_393 = {1{`RANDOM}};
  mem_393 = _RAND_393[18:0];
  _RAND_394 = {1{`RANDOM}};
  mem_394 = _RAND_394[18:0];
  _RAND_395 = {1{`RANDOM}};
  mem_395 = _RAND_395[18:0];
  _RAND_396 = {1{`RANDOM}};
  mem_396 = _RAND_396[18:0];
  _RAND_397 = {1{`RANDOM}};
  mem_397 = _RAND_397[18:0];
  _RAND_398 = {1{`RANDOM}};
  mem_398 = _RAND_398[18:0];
  _RAND_399 = {1{`RANDOM}};
  mem_399 = _RAND_399[18:0];
  _RAND_400 = {1{`RANDOM}};
  mem_400 = _RAND_400[18:0];
  _RAND_401 = {1{`RANDOM}};
  mem_401 = _RAND_401[18:0];
  _RAND_402 = {1{`RANDOM}};
  mem_402 = _RAND_402[18:0];
  _RAND_403 = {1{`RANDOM}};
  mem_403 = _RAND_403[18:0];
  _RAND_404 = {1{`RANDOM}};
  mem_404 = _RAND_404[18:0];
  _RAND_405 = {1{`RANDOM}};
  mem_405 = _RAND_405[18:0];
  _RAND_406 = {1{`RANDOM}};
  mem_406 = _RAND_406[18:0];
  _RAND_407 = {1{`RANDOM}};
  mem_407 = _RAND_407[18:0];
  _RAND_408 = {1{`RANDOM}};
  mem_408 = _RAND_408[18:0];
  _RAND_409 = {1{`RANDOM}};
  mem_409 = _RAND_409[18:0];
  _RAND_410 = {1{`RANDOM}};
  mem_410 = _RAND_410[18:0];
  _RAND_411 = {1{`RANDOM}};
  mem_411 = _RAND_411[18:0];
  _RAND_412 = {1{`RANDOM}};
  mem_412 = _RAND_412[18:0];
  _RAND_413 = {1{`RANDOM}};
  mem_413 = _RAND_413[18:0];
  _RAND_414 = {1{`RANDOM}};
  mem_414 = _RAND_414[18:0];
  _RAND_415 = {1{`RANDOM}};
  mem_415 = _RAND_415[18:0];
  _RAND_416 = {1{`RANDOM}};
  mem_416 = _RAND_416[18:0];
  _RAND_417 = {1{`RANDOM}};
  mem_417 = _RAND_417[18:0];
  _RAND_418 = {1{`RANDOM}};
  mem_418 = _RAND_418[18:0];
  _RAND_419 = {1{`RANDOM}};
  mem_419 = _RAND_419[18:0];
  _RAND_420 = {1{`RANDOM}};
  mem_420 = _RAND_420[18:0];
  _RAND_421 = {1{`RANDOM}};
  mem_421 = _RAND_421[18:0];
  _RAND_422 = {1{`RANDOM}};
  mem_422 = _RAND_422[18:0];
  _RAND_423 = {1{`RANDOM}};
  mem_423 = _RAND_423[18:0];
  _RAND_424 = {1{`RANDOM}};
  mem_424 = _RAND_424[18:0];
  _RAND_425 = {1{`RANDOM}};
  mem_425 = _RAND_425[18:0];
  _RAND_426 = {1{`RANDOM}};
  mem_426 = _RAND_426[18:0];
  _RAND_427 = {1{`RANDOM}};
  mem_427 = _RAND_427[18:0];
  _RAND_428 = {1{`RANDOM}};
  mem_428 = _RAND_428[18:0];
  _RAND_429 = {1{`RANDOM}};
  mem_429 = _RAND_429[18:0];
  _RAND_430 = {1{`RANDOM}};
  mem_430 = _RAND_430[18:0];
  _RAND_431 = {1{`RANDOM}};
  mem_431 = _RAND_431[18:0];
  _RAND_432 = {1{`RANDOM}};
  mem_432 = _RAND_432[18:0];
  _RAND_433 = {1{`RANDOM}};
  mem_433 = _RAND_433[18:0];
  _RAND_434 = {1{`RANDOM}};
  mem_434 = _RAND_434[18:0];
  _RAND_435 = {1{`RANDOM}};
  mem_435 = _RAND_435[18:0];
  _RAND_436 = {1{`RANDOM}};
  mem_436 = _RAND_436[18:0];
  _RAND_437 = {1{`RANDOM}};
  mem_437 = _RAND_437[18:0];
  _RAND_438 = {1{`RANDOM}};
  mem_438 = _RAND_438[18:0];
  _RAND_439 = {1{`RANDOM}};
  mem_439 = _RAND_439[18:0];
  _RAND_440 = {1{`RANDOM}};
  mem_440 = _RAND_440[18:0];
  _RAND_441 = {1{`RANDOM}};
  mem_441 = _RAND_441[18:0];
  _RAND_442 = {1{`RANDOM}};
  mem_442 = _RAND_442[18:0];
  _RAND_443 = {1{`RANDOM}};
  mem_443 = _RAND_443[18:0];
  _RAND_444 = {1{`RANDOM}};
  mem_444 = _RAND_444[18:0];
  _RAND_445 = {1{`RANDOM}};
  mem_445 = _RAND_445[18:0];
  _RAND_446 = {1{`RANDOM}};
  mem_446 = _RAND_446[18:0];
  _RAND_447 = {1{`RANDOM}};
  mem_447 = _RAND_447[18:0];
  _RAND_448 = {1{`RANDOM}};
  mem_448 = _RAND_448[18:0];
  _RAND_449 = {1{`RANDOM}};
  mem_449 = _RAND_449[18:0];
  _RAND_450 = {1{`RANDOM}};
  mem_450 = _RAND_450[18:0];
  _RAND_451 = {1{`RANDOM}};
  mem_451 = _RAND_451[18:0];
  _RAND_452 = {1{`RANDOM}};
  mem_452 = _RAND_452[18:0];
  _RAND_453 = {1{`RANDOM}};
  mem_453 = _RAND_453[18:0];
  _RAND_454 = {1{`RANDOM}};
  mem_454 = _RAND_454[18:0];
  _RAND_455 = {1{`RANDOM}};
  mem_455 = _RAND_455[18:0];
  _RAND_456 = {1{`RANDOM}};
  mem_456 = _RAND_456[18:0];
  _RAND_457 = {1{`RANDOM}};
  mem_457 = _RAND_457[18:0];
  _RAND_458 = {1{`RANDOM}};
  mem_458 = _RAND_458[18:0];
  _RAND_459 = {1{`RANDOM}};
  mem_459 = _RAND_459[18:0];
  _RAND_460 = {1{`RANDOM}};
  mem_460 = _RAND_460[18:0];
  _RAND_461 = {1{`RANDOM}};
  mem_461 = _RAND_461[18:0];
  _RAND_462 = {1{`RANDOM}};
  mem_462 = _RAND_462[18:0];
  _RAND_463 = {1{`RANDOM}};
  mem_463 = _RAND_463[18:0];
  _RAND_464 = {1{`RANDOM}};
  mem_464 = _RAND_464[18:0];
  _RAND_465 = {1{`RANDOM}};
  mem_465 = _RAND_465[18:0];
  _RAND_466 = {1{`RANDOM}};
  mem_466 = _RAND_466[18:0];
  _RAND_467 = {1{`RANDOM}};
  mem_467 = _RAND_467[18:0];
  _RAND_468 = {1{`RANDOM}};
  mem_468 = _RAND_468[18:0];
  _RAND_469 = {1{`RANDOM}};
  mem_469 = _RAND_469[18:0];
  _RAND_470 = {1{`RANDOM}};
  mem_470 = _RAND_470[18:0];
  _RAND_471 = {1{`RANDOM}};
  mem_471 = _RAND_471[18:0];
  _RAND_472 = {1{`RANDOM}};
  mem_472 = _RAND_472[18:0];
  _RAND_473 = {1{`RANDOM}};
  mem_473 = _RAND_473[18:0];
  _RAND_474 = {1{`RANDOM}};
  mem_474 = _RAND_474[18:0];
  _RAND_475 = {1{`RANDOM}};
  mem_475 = _RAND_475[18:0];
  _RAND_476 = {1{`RANDOM}};
  mem_476 = _RAND_476[18:0];
  _RAND_477 = {1{`RANDOM}};
  mem_477 = _RAND_477[18:0];
  _RAND_478 = {1{`RANDOM}};
  mem_478 = _RAND_478[18:0];
  _RAND_479 = {1{`RANDOM}};
  mem_479 = _RAND_479[18:0];
  _RAND_480 = {1{`RANDOM}};
  mem_480 = _RAND_480[18:0];
  _RAND_481 = {1{`RANDOM}};
  mem_481 = _RAND_481[18:0];
  _RAND_482 = {1{`RANDOM}};
  mem_482 = _RAND_482[18:0];
  _RAND_483 = {1{`RANDOM}};
  mem_483 = _RAND_483[18:0];
  _RAND_484 = {1{`RANDOM}};
  mem_484 = _RAND_484[18:0];
  _RAND_485 = {1{`RANDOM}};
  mem_485 = _RAND_485[18:0];
  _RAND_486 = {1{`RANDOM}};
  mem_486 = _RAND_486[18:0];
  _RAND_487 = {1{`RANDOM}};
  mem_487 = _RAND_487[18:0];
  _RAND_488 = {1{`RANDOM}};
  mem_488 = _RAND_488[18:0];
  _RAND_489 = {1{`RANDOM}};
  mem_489 = _RAND_489[18:0];
  _RAND_490 = {1{`RANDOM}};
  mem_490 = _RAND_490[18:0];
  _RAND_491 = {1{`RANDOM}};
  mem_491 = _RAND_491[18:0];
  _RAND_492 = {1{`RANDOM}};
  mem_492 = _RAND_492[18:0];
  _RAND_493 = {1{`RANDOM}};
  mem_493 = _RAND_493[18:0];
  _RAND_494 = {1{`RANDOM}};
  mem_494 = _RAND_494[18:0];
  _RAND_495 = {1{`RANDOM}};
  mem_495 = _RAND_495[18:0];
  _RAND_496 = {1{`RANDOM}};
  mem_496 = _RAND_496[18:0];
  _RAND_497 = {1{`RANDOM}};
  mem_497 = _RAND_497[18:0];
  _RAND_498 = {1{`RANDOM}};
  mem_498 = _RAND_498[18:0];
  _RAND_499 = {1{`RANDOM}};
  mem_499 = _RAND_499[18:0];
  _RAND_500 = {1{`RANDOM}};
  mem_500 = _RAND_500[18:0];
  _RAND_501 = {1{`RANDOM}};
  mem_501 = _RAND_501[18:0];
  _RAND_502 = {1{`RANDOM}};
  mem_502 = _RAND_502[18:0];
  _RAND_503 = {1{`RANDOM}};
  mem_503 = _RAND_503[18:0];
  _RAND_504 = {1{`RANDOM}};
  mem_504 = _RAND_504[18:0];
  _RAND_505 = {1{`RANDOM}};
  mem_505 = _RAND_505[18:0];
  _RAND_506 = {1{`RANDOM}};
  mem_506 = _RAND_506[18:0];
  _RAND_507 = {1{`RANDOM}};
  mem_507 = _RAND_507[18:0];
  _RAND_508 = {1{`RANDOM}};
  mem_508 = _RAND_508[18:0];
  _RAND_509 = {1{`RANDOM}};
  mem_509 = _RAND_509[18:0];
  _RAND_510 = {1{`RANDOM}};
  mem_510 = _RAND_510[18:0];
  _RAND_511 = {1{`RANDOM}};
  mem_511 = _RAND_511[18:0];
  _RAND_512 = {1{`RANDOM}};
  io_dout_REG = _RAND_512[18:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinglePortBRAM_1(
  input         clock,
  input         reset,
  input         io_we,
  input  [8:0]  io_addr,
  input  [18:0] io_din,
  output [18:0] io_dout
);
  wire  sim_single_port_bram_clock; // @[RAMWrapper.scala 275:38]
  wire  sim_single_port_bram_reset; // @[RAMWrapper.scala 275:38]
  wire  sim_single_port_bram_io_we; // @[RAMWrapper.scala 275:38]
  wire [8:0] sim_single_port_bram_io_addr; // @[RAMWrapper.scala 275:38]
  wire [18:0] sim_single_port_bram_io_din; // @[RAMWrapper.scala 275:38]
  wire [18:0] sim_single_port_bram_io_dout; // @[RAMWrapper.scala 275:38]
  SimSinglePortBRAM_1 sim_single_port_bram ( // @[RAMWrapper.scala 275:38]
    .clock(sim_single_port_bram_clock),
    .reset(sim_single_port_bram_reset),
    .io_we(sim_single_port_bram_io_we),
    .io_addr(sim_single_port_bram_io_addr),
    .io_din(sim_single_port_bram_io_din),
    .io_dout(sim_single_port_bram_io_dout)
  );
  assign io_dout = sim_single_port_bram_io_dout; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_clock = clock;
  assign sim_single_port_bram_reset = reset;
  assign sim_single_port_bram_io_we = io_we; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_io_addr = io_addr; // @[RAMWrapper.scala 276:29]
  assign sim_single_port_bram_io_din = io_din; // @[RAMWrapper.scala 276:29]
endmodule
module ICacheMeta(
  input         clock,
  input         reset,
  input         io_we,
  input  [8:0]  io_addr,
  input  [18:0] io_din,
  output [18:0] io_dout
);
  wire  blk_clock; // @[ICache.scala 20:19]
  wire  blk_reset; // @[ICache.scala 20:19]
  wire  blk_io_we; // @[ICache.scala 20:19]
  wire [8:0] blk_io_addr; // @[ICache.scala 20:19]
  wire [18:0] blk_io_din; // @[ICache.scala 20:19]
  wire [18:0] blk_io_dout; // @[ICache.scala 20:19]
  SinglePortBRAM_1 blk ( // @[ICache.scala 20:19]
    .clock(blk_clock),
    .reset(blk_reset),
    .io_we(blk_io_we),
    .io_addr(blk_io_addr),
    .io_din(blk_io_din),
    .io_dout(blk_io_dout)
  );
  assign io_dout = blk_io_dout; // @[ICache.scala 26:16]
  assign blk_clock = clock;
  assign blk_reset = reset;
  assign blk_io_we = io_we; // @[ICache.scala 23:16]
  assign blk_io_addr = io_addr; // @[ICache.scala 24:16]
  assign blk_io_din = io_din; // @[ICache.scala 25:16]
endmodule
module ICache(
  input          clock,
  input          reset,
  input  [31:0]  io_cpu_req_bits_addr,
  input  [2:0]   io_cpu_req_bits_mtype,
  output         io_cpu_resp_valid,
  output [31:0]  io_cpu_resp_bits_rdata_0,
  output [31:0]  io_cpu_resp_bits_rdata_1,
  output         io_cpu_resp_bits_respn,
  output         io_bar_req_valid,
  output [31:0]  io_bar_req_addr,
  input          io_bar_resp_valid,
  input  [255:0] io_bar_resp_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  data_clock; // @[ICache.scala 38:20]
  wire  data_reset; // @[ICache.scala 38:20]
  wire  data_io_we; // @[ICache.scala 38:20]
  wire [8:0] data_io_addr; // @[ICache.scala 38:20]
  wire [255:0] data_io_din; // @[ICache.scala 38:20]
  wire [255:0] data_io_dout; // @[ICache.scala 38:20]
  wire  meta_clock; // @[ICache.scala 39:20]
  wire  meta_reset; // @[ICache.scala 39:20]
  wire  meta_io_we; // @[ICache.scala 39:20]
  wire [8:0] meta_io_addr; // @[ICache.scala 39:20]
  wire [18:0] meta_io_din; // @[ICache.scala 39:20]
  wire [18:0] meta_io_dout; // @[ICache.scala 39:20]
  wire [17:0] tag_req = io_cpu_req_bits_addr[31:14]; // @[ICache.scala 40:39]
  reg [31:0] req_addr; // @[ICache.scala 44:25]
  wire [2:0] word1 = req_addr[4:2]; // @[ICache.scala 45:23]
  wire [2:0] word2 = word1 + 3'h1; // @[ICache.scala 46:21]
  wire  hit = meta_io_dout[18] & meta_io_dout[17:0] == req_addr[31:14]; // @[ICache.scala 48:42]
  reg [31:0] refill_data_0; // @[ICache.scala 55:24]
  reg [31:0] refill_data_1; // @[ICache.scala 55:24]
  reg [31:0] refill_data_2; // @[ICache.scala 55:24]
  reg [31:0] refill_data_3; // @[ICache.scala 55:24]
  reg [31:0] refill_data_4; // @[ICache.scala 55:24]
  reg [31:0] refill_data_5; // @[ICache.scala 55:24]
  reg [31:0] refill_data_6; // @[ICache.scala 55:24]
  reg [31:0] refill_data_7; // @[ICache.scala 55:24]
  wire [31:0] line_0 = data_io_dout[31:0]; // @[ICache.scala 63:28]
  wire [31:0] line_1 = data_io_dout[63:32]; // @[ICache.scala 63:28]
  wire [31:0] line_2 = data_io_dout[95:64]; // @[ICache.scala 63:28]
  wire [31:0] line_3 = data_io_dout[127:96]; // @[ICache.scala 63:28]
  wire [31:0] line_4 = data_io_dout[159:128]; // @[ICache.scala 63:28]
  wire [31:0] line_5 = data_io_dout[191:160]; // @[ICache.scala 63:28]
  wire [31:0] line_6 = data_io_dout[223:192]; // @[ICache.scala 63:28]
  wire [31:0] line_7 = data_io_dout[255:224]; // @[ICache.scala 63:28]
  reg [1:0] state; // @[ICache.scala 68:22]
  wire  _io_cpu_resp_valid_T = state == 2'h3; // @[ICache.scala 75:30]
  wire [2:0] _io_cpu_resp_bits_respn_T_3 = io_cpu_req_bits_addr[4:2] + 3'h1; // @[ICache.scala 77:47]
  wire  _io_cpu_resp_bits_respn_T_4 = _io_cpu_resp_bits_respn_T_3 != 3'h0; // @[ICache.scala 77:53]
  wire [31:0] _GEN_1 = 3'h1 == word1 ? refill_data_1 : refill_data_0; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_2 = 3'h2 == word1 ? refill_data_2 : _GEN_1; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_3 = 3'h3 == word1 ? refill_data_3 : _GEN_2; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_4 = 3'h4 == word1 ? refill_data_4 : _GEN_3; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_5 = 3'h5 == word1 ? refill_data_5 : _GEN_4; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_6 = 3'h6 == word1 ? refill_data_6 : _GEN_5; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_7 = 3'h7 == word1 ? refill_data_7 : _GEN_6; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_9 = 3'h1 == word1 ? line_1 : line_0; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_10 = 3'h2 == word1 ? line_2 : _GEN_9; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_11 = 3'h3 == word1 ? line_3 : _GEN_10; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_12 = 3'h4 == word1 ? line_4 : _GEN_11; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_13 = 3'h5 == word1 ? line_5 : _GEN_12; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_14 = 3'h6 == word1 ? line_6 : _GEN_13; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_15 = 3'h7 == word1 ? line_7 : _GEN_14; // @[ICache.scala 78:35 ICache.scala 78:35]
  wire [31:0] _GEN_17 = 3'h1 == word2 ? refill_data_1 : refill_data_0; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_18 = 3'h2 == word2 ? refill_data_2 : _GEN_17; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_19 = 3'h3 == word2 ? refill_data_3 : _GEN_18; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_20 = 3'h4 == word2 ? refill_data_4 : _GEN_19; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_21 = 3'h5 == word2 ? refill_data_5 : _GEN_20; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_22 = 3'h6 == word2 ? refill_data_6 : _GEN_21; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_23 = 3'h7 == word2 ? refill_data_7 : _GEN_22; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_25 = 3'h1 == word2 ? line_1 : line_0; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_26 = 3'h2 == word2 ? line_2 : _GEN_25; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_27 = 3'h3 == word2 ? line_3 : _GEN_26; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_28 = 3'h4 == word2 ? line_4 : _GEN_27; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_29 = 3'h5 == word2 ? line_5 : _GEN_28; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_30 = 3'h6 == word2 ? line_6 : _GEN_29; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [31:0] _GEN_31 = 3'h7 == word2 ? line_7 : _GEN_30; // @[ICache.scala 79:35 ICache.scala 79:35]
  wire [26:0] io_bar_req_addr_hi = req_addr[31:5]; // @[ICache.scala 90:13]
  wire [31:0] _io_bar_req_addr_T = {io_bar_req_addr_hi,5'h0}; // @[Cat.scala 30:58]
  wire  _T_1 = ~hit; // @[ICache.scala 104:13]
  wire  _io_bar_req_valid_T = ~io_bar_resp_valid; // @[ICache.scala 111:27]
  wire [1:0] _GEN_34 = io_bar_resp_valid ? 2'h3 : state; // @[ICache.scala 116:30 ICache.scala 121:16]
  wire [29:0] io_bar_req_addr_hi_1 = req_addr[31:2]; // @[ICache.scala 130:36]
  wire [31:0] _io_bar_req_addr_T_1 = {io_bar_req_addr_hi_1,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _io_bar_req_addr_T_3 = _io_bar_req_addr_T_1 + 32'h4; // @[ICache.scala 130:61]
  wire [31:0] _GEN_44 = state == 2'h2 ? _io_bar_req_addr_T_3 : _io_bar_req_addr_T; // @[ICache.scala 129:41 ICache.scala 130:21 ICache.scala 89:19]
  wire  _GEN_45 = state == 2'h2 & _io_bar_req_valid_T; // @[ICache.scala 129:41 ICache.scala 131:22 ICache.scala 87:20]
  wire  _GEN_47 = state == 2'h1 ? ~io_bar_resp_valid : _GEN_45; // @[ICache.scala 109:34 ICache.scala 111:24]
  wire  _GEN_57 = state == 2'h1 & io_bar_resp_valid; // @[ICache.scala 109:34 ICache.scala 49:16]
  wire [31:0] _GEN_58 = state == 2'h1 ? _io_bar_req_addr_T : _GEN_44; // @[ICache.scala 109:34 ICache.scala 89:19]
  SinglePortBRAM data ( // @[ICache.scala 38:20]
    .clock(data_clock),
    .reset(data_reset),
    .io_we(data_io_we),
    .io_addr(data_io_addr),
    .io_din(data_io_din),
    .io_dout(data_io_dout)
  );
  ICacheMeta meta ( // @[ICache.scala 39:20]
    .clock(meta_clock),
    .reset(meta_reset),
    .io_we(meta_io_we),
    .io_addr(meta_io_addr),
    .io_din(meta_io_din),
    .io_dout(meta_io_dout)
  );
  assign io_cpu_resp_valid = state == 2'h3 | hit; // @[ICache.scala 75:43]
  assign io_cpu_resp_bits_rdata_0 = _io_cpu_resp_valid_T ? _GEN_7 : _GEN_15; // @[ICache.scala 78:35]
  assign io_cpu_resp_bits_rdata_1 = _io_cpu_resp_valid_T ? _GEN_23 : _GEN_31; // @[ICache.scala 79:35]
  assign io_cpu_resp_bits_respn = io_cpu_req_bits_mtype == 3'h3 & _io_cpu_resp_bits_respn_T_4; // @[ICache.scala 76:68]
  assign io_bar_req_valid = state == 2'h0 ? _T_1 : _GEN_47; // @[ICache.scala 99:29]
  assign io_bar_req_addr = state == 2'h0 ? _io_bar_req_addr_T : _GEN_58; // @[ICache.scala 99:29 ICache.scala 89:19]
  assign data_clock = clock;
  assign data_reset = reset;
  assign data_io_we = state == 2'h0 ? 1'h0 : _GEN_57; // @[ICache.scala 99:29 ICache.scala 49:16]
  assign data_io_addr = io_cpu_req_bits_addr[13:5]; // @[ICache.scala 41:39]
  assign data_io_din = io_bar_resp_data; // @[ICache.scala 60:15]
  assign meta_clock = clock;
  assign meta_reset = reset;
  assign meta_io_we = state == 2'h0 ? 1'h0 : _GEN_57; // @[ICache.scala 99:29 ICache.scala 49:16]
  assign meta_io_addr = io_cpu_req_bits_addr[13:5]; // @[ICache.scala 41:39]
  assign meta_io_din = {1'h1,tag_req}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    req_addr <= io_cpu_req_bits_addr; // @[ICache.scala 44:25]
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_0 <= io_bar_resp_data[31:0]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_1 <= io_bar_resp_data[63:32]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_2 <= io_bar_resp_data[95:64]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_3 <= io_bar_resp_data[127:96]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_4 <= io_bar_resp_data[159:128]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_5 <= io_bar_resp_data[191:160]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_6 <= io_bar_resp_data[223:192]; // @[ICache.scala 123:26]
        end
      end
    end
    if (!(state == 2'h0)) begin // @[ICache.scala 99:29]
      if (state == 2'h1) begin // @[ICache.scala 109:34]
        if (io_bar_resp_valid) begin // @[ICache.scala 116:30]
          refill_data_7 <= io_bar_resp_data[255:224]; // @[ICache.scala 123:26]
        end
      end
    end
    if (reset) begin // @[ICache.scala 68:22]
      state <= 2'h0; // @[ICache.scala 68:22]
    end else if (state == 2'h0) begin // @[ICache.scala 99:29]
      if (~hit) begin // @[ICache.scala 104:19]
        state <= 2'h1; // @[ICache.scala 105:16]
      end
    end else if (state == 2'h1) begin // @[ICache.scala 109:34]
      state <= _GEN_34;
    end else if (state == 2'h2) begin // @[ICache.scala 129:41]
      state <= _GEN_34; // @[ICache.scala 132:12]
    end else begin
      state <= 2'h0; // @[ICache.scala 134:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  req_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  refill_data_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  refill_data_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  refill_data_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  refill_data_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  refill_data_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  refill_data_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  refill_data_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  refill_data_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimDualPortBRAM_2(
  input          clock,
  input          reset,
  input          io_web,
  input  [8:0]   io_addra,
  input  [8:0]   io_addrb,
  input  [255:0] io_dinb,
  output [255:0] io_douta
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [255:0] _RAND_2;
  reg [255:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [255:0] _RAND_5;
  reg [255:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [255:0] _RAND_9;
  reg [255:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [255:0] _RAND_12;
  reg [255:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [255:0] _RAND_16;
  reg [255:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [255:0] _RAND_22;
  reg [255:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [255:0] _RAND_26;
  reg [255:0] _RAND_27;
  reg [255:0] _RAND_28;
  reg [255:0] _RAND_29;
  reg [255:0] _RAND_30;
  reg [255:0] _RAND_31;
  reg [255:0] _RAND_32;
  reg [255:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [255:0] _RAND_35;
  reg [255:0] _RAND_36;
  reg [255:0] _RAND_37;
  reg [255:0] _RAND_38;
  reg [255:0] _RAND_39;
  reg [255:0] _RAND_40;
  reg [255:0] _RAND_41;
  reg [255:0] _RAND_42;
  reg [255:0] _RAND_43;
  reg [255:0] _RAND_44;
  reg [255:0] _RAND_45;
  reg [255:0] _RAND_46;
  reg [255:0] _RAND_47;
  reg [255:0] _RAND_48;
  reg [255:0] _RAND_49;
  reg [255:0] _RAND_50;
  reg [255:0] _RAND_51;
  reg [255:0] _RAND_52;
  reg [255:0] _RAND_53;
  reg [255:0] _RAND_54;
  reg [255:0] _RAND_55;
  reg [255:0] _RAND_56;
  reg [255:0] _RAND_57;
  reg [255:0] _RAND_58;
  reg [255:0] _RAND_59;
  reg [255:0] _RAND_60;
  reg [255:0] _RAND_61;
  reg [255:0] _RAND_62;
  reg [255:0] _RAND_63;
  reg [255:0] _RAND_64;
  reg [255:0] _RAND_65;
  reg [255:0] _RAND_66;
  reg [255:0] _RAND_67;
  reg [255:0] _RAND_68;
  reg [255:0] _RAND_69;
  reg [255:0] _RAND_70;
  reg [255:0] _RAND_71;
  reg [255:0] _RAND_72;
  reg [255:0] _RAND_73;
  reg [255:0] _RAND_74;
  reg [255:0] _RAND_75;
  reg [255:0] _RAND_76;
  reg [255:0] _RAND_77;
  reg [255:0] _RAND_78;
  reg [255:0] _RAND_79;
  reg [255:0] _RAND_80;
  reg [255:0] _RAND_81;
  reg [255:0] _RAND_82;
  reg [255:0] _RAND_83;
  reg [255:0] _RAND_84;
  reg [255:0] _RAND_85;
  reg [255:0] _RAND_86;
  reg [255:0] _RAND_87;
  reg [255:0] _RAND_88;
  reg [255:0] _RAND_89;
  reg [255:0] _RAND_90;
  reg [255:0] _RAND_91;
  reg [255:0] _RAND_92;
  reg [255:0] _RAND_93;
  reg [255:0] _RAND_94;
  reg [255:0] _RAND_95;
  reg [255:0] _RAND_96;
  reg [255:0] _RAND_97;
  reg [255:0] _RAND_98;
  reg [255:0] _RAND_99;
  reg [255:0] _RAND_100;
  reg [255:0] _RAND_101;
  reg [255:0] _RAND_102;
  reg [255:0] _RAND_103;
  reg [255:0] _RAND_104;
  reg [255:0] _RAND_105;
  reg [255:0] _RAND_106;
  reg [255:0] _RAND_107;
  reg [255:0] _RAND_108;
  reg [255:0] _RAND_109;
  reg [255:0] _RAND_110;
  reg [255:0] _RAND_111;
  reg [255:0] _RAND_112;
  reg [255:0] _RAND_113;
  reg [255:0] _RAND_114;
  reg [255:0] _RAND_115;
  reg [255:0] _RAND_116;
  reg [255:0] _RAND_117;
  reg [255:0] _RAND_118;
  reg [255:0] _RAND_119;
  reg [255:0] _RAND_120;
  reg [255:0] _RAND_121;
  reg [255:0] _RAND_122;
  reg [255:0] _RAND_123;
  reg [255:0] _RAND_124;
  reg [255:0] _RAND_125;
  reg [255:0] _RAND_126;
  reg [255:0] _RAND_127;
  reg [255:0] _RAND_128;
  reg [255:0] _RAND_129;
  reg [255:0] _RAND_130;
  reg [255:0] _RAND_131;
  reg [255:0] _RAND_132;
  reg [255:0] _RAND_133;
  reg [255:0] _RAND_134;
  reg [255:0] _RAND_135;
  reg [255:0] _RAND_136;
  reg [255:0] _RAND_137;
  reg [255:0] _RAND_138;
  reg [255:0] _RAND_139;
  reg [255:0] _RAND_140;
  reg [255:0] _RAND_141;
  reg [255:0] _RAND_142;
  reg [255:0] _RAND_143;
  reg [255:0] _RAND_144;
  reg [255:0] _RAND_145;
  reg [255:0] _RAND_146;
  reg [255:0] _RAND_147;
  reg [255:0] _RAND_148;
  reg [255:0] _RAND_149;
  reg [255:0] _RAND_150;
  reg [255:0] _RAND_151;
  reg [255:0] _RAND_152;
  reg [255:0] _RAND_153;
  reg [255:0] _RAND_154;
  reg [255:0] _RAND_155;
  reg [255:0] _RAND_156;
  reg [255:0] _RAND_157;
  reg [255:0] _RAND_158;
  reg [255:0] _RAND_159;
  reg [255:0] _RAND_160;
  reg [255:0] _RAND_161;
  reg [255:0] _RAND_162;
  reg [255:0] _RAND_163;
  reg [255:0] _RAND_164;
  reg [255:0] _RAND_165;
  reg [255:0] _RAND_166;
  reg [255:0] _RAND_167;
  reg [255:0] _RAND_168;
  reg [255:0] _RAND_169;
  reg [255:0] _RAND_170;
  reg [255:0] _RAND_171;
  reg [255:0] _RAND_172;
  reg [255:0] _RAND_173;
  reg [255:0] _RAND_174;
  reg [255:0] _RAND_175;
  reg [255:0] _RAND_176;
  reg [255:0] _RAND_177;
  reg [255:0] _RAND_178;
  reg [255:0] _RAND_179;
  reg [255:0] _RAND_180;
  reg [255:0] _RAND_181;
  reg [255:0] _RAND_182;
  reg [255:0] _RAND_183;
  reg [255:0] _RAND_184;
  reg [255:0] _RAND_185;
  reg [255:0] _RAND_186;
  reg [255:0] _RAND_187;
  reg [255:0] _RAND_188;
  reg [255:0] _RAND_189;
  reg [255:0] _RAND_190;
  reg [255:0] _RAND_191;
  reg [255:0] _RAND_192;
  reg [255:0] _RAND_193;
  reg [255:0] _RAND_194;
  reg [255:0] _RAND_195;
  reg [255:0] _RAND_196;
  reg [255:0] _RAND_197;
  reg [255:0] _RAND_198;
  reg [255:0] _RAND_199;
  reg [255:0] _RAND_200;
  reg [255:0] _RAND_201;
  reg [255:0] _RAND_202;
  reg [255:0] _RAND_203;
  reg [255:0] _RAND_204;
  reg [255:0] _RAND_205;
  reg [255:0] _RAND_206;
  reg [255:0] _RAND_207;
  reg [255:0] _RAND_208;
  reg [255:0] _RAND_209;
  reg [255:0] _RAND_210;
  reg [255:0] _RAND_211;
  reg [255:0] _RAND_212;
  reg [255:0] _RAND_213;
  reg [255:0] _RAND_214;
  reg [255:0] _RAND_215;
  reg [255:0] _RAND_216;
  reg [255:0] _RAND_217;
  reg [255:0] _RAND_218;
  reg [255:0] _RAND_219;
  reg [255:0] _RAND_220;
  reg [255:0] _RAND_221;
  reg [255:0] _RAND_222;
  reg [255:0] _RAND_223;
  reg [255:0] _RAND_224;
  reg [255:0] _RAND_225;
  reg [255:0] _RAND_226;
  reg [255:0] _RAND_227;
  reg [255:0] _RAND_228;
  reg [255:0] _RAND_229;
  reg [255:0] _RAND_230;
  reg [255:0] _RAND_231;
  reg [255:0] _RAND_232;
  reg [255:0] _RAND_233;
  reg [255:0] _RAND_234;
  reg [255:0] _RAND_235;
  reg [255:0] _RAND_236;
  reg [255:0] _RAND_237;
  reg [255:0] _RAND_238;
  reg [255:0] _RAND_239;
  reg [255:0] _RAND_240;
  reg [255:0] _RAND_241;
  reg [255:0] _RAND_242;
  reg [255:0] _RAND_243;
  reg [255:0] _RAND_244;
  reg [255:0] _RAND_245;
  reg [255:0] _RAND_246;
  reg [255:0] _RAND_247;
  reg [255:0] _RAND_248;
  reg [255:0] _RAND_249;
  reg [255:0] _RAND_250;
  reg [255:0] _RAND_251;
  reg [255:0] _RAND_252;
  reg [255:0] _RAND_253;
  reg [255:0] _RAND_254;
  reg [255:0] _RAND_255;
  reg [255:0] _RAND_256;
  reg [255:0] _RAND_257;
  reg [255:0] _RAND_258;
  reg [255:0] _RAND_259;
  reg [255:0] _RAND_260;
  reg [255:0] _RAND_261;
  reg [255:0] _RAND_262;
  reg [255:0] _RAND_263;
  reg [255:0] _RAND_264;
  reg [255:0] _RAND_265;
  reg [255:0] _RAND_266;
  reg [255:0] _RAND_267;
  reg [255:0] _RAND_268;
  reg [255:0] _RAND_269;
  reg [255:0] _RAND_270;
  reg [255:0] _RAND_271;
  reg [255:0] _RAND_272;
  reg [255:0] _RAND_273;
  reg [255:0] _RAND_274;
  reg [255:0] _RAND_275;
  reg [255:0] _RAND_276;
  reg [255:0] _RAND_277;
  reg [255:0] _RAND_278;
  reg [255:0] _RAND_279;
  reg [255:0] _RAND_280;
  reg [255:0] _RAND_281;
  reg [255:0] _RAND_282;
  reg [255:0] _RAND_283;
  reg [255:0] _RAND_284;
  reg [255:0] _RAND_285;
  reg [255:0] _RAND_286;
  reg [255:0] _RAND_287;
  reg [255:0] _RAND_288;
  reg [255:0] _RAND_289;
  reg [255:0] _RAND_290;
  reg [255:0] _RAND_291;
  reg [255:0] _RAND_292;
  reg [255:0] _RAND_293;
  reg [255:0] _RAND_294;
  reg [255:0] _RAND_295;
  reg [255:0] _RAND_296;
  reg [255:0] _RAND_297;
  reg [255:0] _RAND_298;
  reg [255:0] _RAND_299;
  reg [255:0] _RAND_300;
  reg [255:0] _RAND_301;
  reg [255:0] _RAND_302;
  reg [255:0] _RAND_303;
  reg [255:0] _RAND_304;
  reg [255:0] _RAND_305;
  reg [255:0] _RAND_306;
  reg [255:0] _RAND_307;
  reg [255:0] _RAND_308;
  reg [255:0] _RAND_309;
  reg [255:0] _RAND_310;
  reg [255:0] _RAND_311;
  reg [255:0] _RAND_312;
  reg [255:0] _RAND_313;
  reg [255:0] _RAND_314;
  reg [255:0] _RAND_315;
  reg [255:0] _RAND_316;
  reg [255:0] _RAND_317;
  reg [255:0] _RAND_318;
  reg [255:0] _RAND_319;
  reg [255:0] _RAND_320;
  reg [255:0] _RAND_321;
  reg [255:0] _RAND_322;
  reg [255:0] _RAND_323;
  reg [255:0] _RAND_324;
  reg [255:0] _RAND_325;
  reg [255:0] _RAND_326;
  reg [255:0] _RAND_327;
  reg [255:0] _RAND_328;
  reg [255:0] _RAND_329;
  reg [255:0] _RAND_330;
  reg [255:0] _RAND_331;
  reg [255:0] _RAND_332;
  reg [255:0] _RAND_333;
  reg [255:0] _RAND_334;
  reg [255:0] _RAND_335;
  reg [255:0] _RAND_336;
  reg [255:0] _RAND_337;
  reg [255:0] _RAND_338;
  reg [255:0] _RAND_339;
  reg [255:0] _RAND_340;
  reg [255:0] _RAND_341;
  reg [255:0] _RAND_342;
  reg [255:0] _RAND_343;
  reg [255:0] _RAND_344;
  reg [255:0] _RAND_345;
  reg [255:0] _RAND_346;
  reg [255:0] _RAND_347;
  reg [255:0] _RAND_348;
  reg [255:0] _RAND_349;
  reg [255:0] _RAND_350;
  reg [255:0] _RAND_351;
  reg [255:0] _RAND_352;
  reg [255:0] _RAND_353;
  reg [255:0] _RAND_354;
  reg [255:0] _RAND_355;
  reg [255:0] _RAND_356;
  reg [255:0] _RAND_357;
  reg [255:0] _RAND_358;
  reg [255:0] _RAND_359;
  reg [255:0] _RAND_360;
  reg [255:0] _RAND_361;
  reg [255:0] _RAND_362;
  reg [255:0] _RAND_363;
  reg [255:0] _RAND_364;
  reg [255:0] _RAND_365;
  reg [255:0] _RAND_366;
  reg [255:0] _RAND_367;
  reg [255:0] _RAND_368;
  reg [255:0] _RAND_369;
  reg [255:0] _RAND_370;
  reg [255:0] _RAND_371;
  reg [255:0] _RAND_372;
  reg [255:0] _RAND_373;
  reg [255:0] _RAND_374;
  reg [255:0] _RAND_375;
  reg [255:0] _RAND_376;
  reg [255:0] _RAND_377;
  reg [255:0] _RAND_378;
  reg [255:0] _RAND_379;
  reg [255:0] _RAND_380;
  reg [255:0] _RAND_381;
  reg [255:0] _RAND_382;
  reg [255:0] _RAND_383;
  reg [255:0] _RAND_384;
  reg [255:0] _RAND_385;
  reg [255:0] _RAND_386;
  reg [255:0] _RAND_387;
  reg [255:0] _RAND_388;
  reg [255:0] _RAND_389;
  reg [255:0] _RAND_390;
  reg [255:0] _RAND_391;
  reg [255:0] _RAND_392;
  reg [255:0] _RAND_393;
  reg [255:0] _RAND_394;
  reg [255:0] _RAND_395;
  reg [255:0] _RAND_396;
  reg [255:0] _RAND_397;
  reg [255:0] _RAND_398;
  reg [255:0] _RAND_399;
  reg [255:0] _RAND_400;
  reg [255:0] _RAND_401;
  reg [255:0] _RAND_402;
  reg [255:0] _RAND_403;
  reg [255:0] _RAND_404;
  reg [255:0] _RAND_405;
  reg [255:0] _RAND_406;
  reg [255:0] _RAND_407;
  reg [255:0] _RAND_408;
  reg [255:0] _RAND_409;
  reg [255:0] _RAND_410;
  reg [255:0] _RAND_411;
  reg [255:0] _RAND_412;
  reg [255:0] _RAND_413;
  reg [255:0] _RAND_414;
  reg [255:0] _RAND_415;
  reg [255:0] _RAND_416;
  reg [255:0] _RAND_417;
  reg [255:0] _RAND_418;
  reg [255:0] _RAND_419;
  reg [255:0] _RAND_420;
  reg [255:0] _RAND_421;
  reg [255:0] _RAND_422;
  reg [255:0] _RAND_423;
  reg [255:0] _RAND_424;
  reg [255:0] _RAND_425;
  reg [255:0] _RAND_426;
  reg [255:0] _RAND_427;
  reg [255:0] _RAND_428;
  reg [255:0] _RAND_429;
  reg [255:0] _RAND_430;
  reg [255:0] _RAND_431;
  reg [255:0] _RAND_432;
  reg [255:0] _RAND_433;
  reg [255:0] _RAND_434;
  reg [255:0] _RAND_435;
  reg [255:0] _RAND_436;
  reg [255:0] _RAND_437;
  reg [255:0] _RAND_438;
  reg [255:0] _RAND_439;
  reg [255:0] _RAND_440;
  reg [255:0] _RAND_441;
  reg [255:0] _RAND_442;
  reg [255:0] _RAND_443;
  reg [255:0] _RAND_444;
  reg [255:0] _RAND_445;
  reg [255:0] _RAND_446;
  reg [255:0] _RAND_447;
  reg [255:0] _RAND_448;
  reg [255:0] _RAND_449;
  reg [255:0] _RAND_450;
  reg [255:0] _RAND_451;
  reg [255:0] _RAND_452;
  reg [255:0] _RAND_453;
  reg [255:0] _RAND_454;
  reg [255:0] _RAND_455;
  reg [255:0] _RAND_456;
  reg [255:0] _RAND_457;
  reg [255:0] _RAND_458;
  reg [255:0] _RAND_459;
  reg [255:0] _RAND_460;
  reg [255:0] _RAND_461;
  reg [255:0] _RAND_462;
  reg [255:0] _RAND_463;
  reg [255:0] _RAND_464;
  reg [255:0] _RAND_465;
  reg [255:0] _RAND_466;
  reg [255:0] _RAND_467;
  reg [255:0] _RAND_468;
  reg [255:0] _RAND_469;
  reg [255:0] _RAND_470;
  reg [255:0] _RAND_471;
  reg [255:0] _RAND_472;
  reg [255:0] _RAND_473;
  reg [255:0] _RAND_474;
  reg [255:0] _RAND_475;
  reg [255:0] _RAND_476;
  reg [255:0] _RAND_477;
  reg [255:0] _RAND_478;
  reg [255:0] _RAND_479;
  reg [255:0] _RAND_480;
  reg [255:0] _RAND_481;
  reg [255:0] _RAND_482;
  reg [255:0] _RAND_483;
  reg [255:0] _RAND_484;
  reg [255:0] _RAND_485;
  reg [255:0] _RAND_486;
  reg [255:0] _RAND_487;
  reg [255:0] _RAND_488;
  reg [255:0] _RAND_489;
  reg [255:0] _RAND_490;
  reg [255:0] _RAND_491;
  reg [255:0] _RAND_492;
  reg [255:0] _RAND_493;
  reg [255:0] _RAND_494;
  reg [255:0] _RAND_495;
  reg [255:0] _RAND_496;
  reg [255:0] _RAND_497;
  reg [255:0] _RAND_498;
  reg [255:0] _RAND_499;
  reg [255:0] _RAND_500;
  reg [255:0] _RAND_501;
  reg [255:0] _RAND_502;
  reg [255:0] _RAND_503;
  reg [255:0] _RAND_504;
  reg [255:0] _RAND_505;
  reg [255:0] _RAND_506;
  reg [255:0] _RAND_507;
  reg [255:0] _RAND_508;
  reg [255:0] _RAND_509;
  reg [255:0] _RAND_510;
  reg [255:0] _RAND_511;
  reg [255:0] _RAND_512;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] mem_0; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_1; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_2; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_3; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_4; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_5; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_6; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_7; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_8; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_9; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_10; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_11; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_12; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_13; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_14; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_15; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_16; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_17; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_18; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_19; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_20; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_21; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_22; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_23; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_24; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_25; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_26; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_27; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_28; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_29; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_30; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_31; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_32; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_33; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_34; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_35; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_36; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_37; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_38; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_39; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_40; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_41; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_42; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_43; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_44; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_45; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_46; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_47; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_48; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_49; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_50; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_51; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_52; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_53; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_54; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_55; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_56; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_57; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_58; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_59; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_60; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_61; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_62; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_63; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_64; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_65; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_66; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_67; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_68; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_69; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_70; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_71; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_72; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_73; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_74; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_75; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_76; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_77; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_78; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_79; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_80; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_81; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_82; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_83; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_84; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_85; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_86; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_87; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_88; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_89; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_90; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_91; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_92; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_93; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_94; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_95; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_96; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_97; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_98; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_99; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_100; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_101; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_102; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_103; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_104; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_105; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_106; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_107; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_108; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_109; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_110; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_111; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_112; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_113; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_114; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_115; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_116; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_117; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_118; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_119; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_120; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_121; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_122; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_123; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_124; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_125; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_126; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_127; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_128; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_129; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_130; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_131; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_132; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_133; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_134; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_135; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_136; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_137; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_138; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_139; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_140; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_141; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_142; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_143; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_144; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_145; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_146; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_147; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_148; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_149; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_150; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_151; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_152; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_153; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_154; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_155; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_156; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_157; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_158; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_159; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_160; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_161; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_162; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_163; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_164; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_165; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_166; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_167; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_168; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_169; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_170; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_171; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_172; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_173; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_174; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_175; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_176; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_177; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_178; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_179; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_180; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_181; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_182; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_183; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_184; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_185; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_186; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_187; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_188; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_189; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_190; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_191; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_192; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_193; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_194; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_195; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_196; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_197; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_198; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_199; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_200; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_201; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_202; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_203; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_204; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_205; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_206; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_207; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_208; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_209; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_210; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_211; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_212; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_213; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_214; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_215; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_216; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_217; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_218; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_219; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_220; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_221; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_222; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_223; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_224; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_225; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_226; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_227; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_228; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_229; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_230; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_231; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_232; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_233; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_234; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_235; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_236; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_237; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_238; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_239; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_240; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_241; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_242; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_243; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_244; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_245; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_246; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_247; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_248; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_249; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_250; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_251; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_252; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_253; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_254; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_255; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_256; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_257; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_258; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_259; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_260; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_261; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_262; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_263; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_264; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_265; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_266; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_267; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_268; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_269; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_270; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_271; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_272; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_273; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_274; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_275; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_276; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_277; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_278; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_279; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_280; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_281; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_282; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_283; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_284; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_285; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_286; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_287; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_288; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_289; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_290; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_291; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_292; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_293; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_294; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_295; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_296; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_297; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_298; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_299; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_300; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_301; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_302; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_303; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_304; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_305; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_306; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_307; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_308; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_309; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_310; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_311; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_312; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_313; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_314; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_315; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_316; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_317; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_318; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_319; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_320; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_321; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_322; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_323; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_324; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_325; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_326; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_327; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_328; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_329; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_330; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_331; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_332; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_333; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_334; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_335; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_336; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_337; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_338; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_339; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_340; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_341; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_342; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_343; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_344; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_345; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_346; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_347; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_348; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_349; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_350; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_351; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_352; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_353; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_354; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_355; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_356; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_357; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_358; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_359; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_360; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_361; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_362; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_363; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_364; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_365; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_366; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_367; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_368; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_369; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_370; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_371; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_372; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_373; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_374; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_375; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_376; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_377; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_378; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_379; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_380; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_381; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_382; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_383; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_384; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_385; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_386; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_387; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_388; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_389; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_390; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_391; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_392; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_393; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_394; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_395; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_396; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_397; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_398; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_399; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_400; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_401; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_402; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_403; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_404; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_405; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_406; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_407; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_408; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_409; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_410; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_411; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_412; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_413; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_414; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_415; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_416; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_417; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_418; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_419; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_420; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_421; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_422; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_423; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_424; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_425; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_426; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_427; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_428; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_429; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_430; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_431; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_432; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_433; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_434; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_435; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_436; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_437; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_438; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_439; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_440; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_441; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_442; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_443; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_444; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_445; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_446; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_447; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_448; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_449; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_450; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_451; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_452; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_453; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_454; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_455; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_456; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_457; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_458; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_459; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_460; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_461; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_462; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_463; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_464; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_465; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_466; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_467; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_468; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_469; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_470; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_471; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_472; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_473; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_474; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_475; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_476; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_477; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_478; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_479; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_480; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_481; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_482; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_483; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_484; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_485; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_486; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_487; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_488; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_489; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_490; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_491; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_492; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_493; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_494; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_495; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_496; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_497; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_498; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_499; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_500; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_501; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_502; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_503; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_504; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_505; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_506; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_507; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_508; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_509; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_510; // @[RAMWrapper.scala 41:20]
  reg [255:0] mem_511; // @[RAMWrapper.scala 41:20]
  reg [255:0] io_douta_REG; // @[RAMWrapper.scala 43:22]
  wire [255:0] _GEN_1 = 9'h1 == io_addra ? mem_1 : mem_0; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_2 = 9'h2 == io_addra ? mem_2 : _GEN_1; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_3 = 9'h3 == io_addra ? mem_3 : _GEN_2; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_4 = 9'h4 == io_addra ? mem_4 : _GEN_3; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_5 = 9'h5 == io_addra ? mem_5 : _GEN_4; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_6 = 9'h6 == io_addra ? mem_6 : _GEN_5; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_7 = 9'h7 == io_addra ? mem_7 : _GEN_6; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_8 = 9'h8 == io_addra ? mem_8 : _GEN_7; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_9 = 9'h9 == io_addra ? mem_9 : _GEN_8; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_10 = 9'ha == io_addra ? mem_10 : _GEN_9; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_11 = 9'hb == io_addra ? mem_11 : _GEN_10; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_12 = 9'hc == io_addra ? mem_12 : _GEN_11; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_13 = 9'hd == io_addra ? mem_13 : _GEN_12; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_14 = 9'he == io_addra ? mem_14 : _GEN_13; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_15 = 9'hf == io_addra ? mem_15 : _GEN_14; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_16 = 9'h10 == io_addra ? mem_16 : _GEN_15; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_17 = 9'h11 == io_addra ? mem_17 : _GEN_16; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_18 = 9'h12 == io_addra ? mem_18 : _GEN_17; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_19 = 9'h13 == io_addra ? mem_19 : _GEN_18; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_20 = 9'h14 == io_addra ? mem_20 : _GEN_19; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_21 = 9'h15 == io_addra ? mem_21 : _GEN_20; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_22 = 9'h16 == io_addra ? mem_22 : _GEN_21; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_23 = 9'h17 == io_addra ? mem_23 : _GEN_22; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_24 = 9'h18 == io_addra ? mem_24 : _GEN_23; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_25 = 9'h19 == io_addra ? mem_25 : _GEN_24; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_26 = 9'h1a == io_addra ? mem_26 : _GEN_25; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_27 = 9'h1b == io_addra ? mem_27 : _GEN_26; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_28 = 9'h1c == io_addra ? mem_28 : _GEN_27; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_29 = 9'h1d == io_addra ? mem_29 : _GEN_28; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_30 = 9'h1e == io_addra ? mem_30 : _GEN_29; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_31 = 9'h1f == io_addra ? mem_31 : _GEN_30; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_32 = 9'h20 == io_addra ? mem_32 : _GEN_31; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_33 = 9'h21 == io_addra ? mem_33 : _GEN_32; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_34 = 9'h22 == io_addra ? mem_34 : _GEN_33; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_35 = 9'h23 == io_addra ? mem_35 : _GEN_34; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_36 = 9'h24 == io_addra ? mem_36 : _GEN_35; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_37 = 9'h25 == io_addra ? mem_37 : _GEN_36; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_38 = 9'h26 == io_addra ? mem_38 : _GEN_37; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_39 = 9'h27 == io_addra ? mem_39 : _GEN_38; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_40 = 9'h28 == io_addra ? mem_40 : _GEN_39; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_41 = 9'h29 == io_addra ? mem_41 : _GEN_40; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_42 = 9'h2a == io_addra ? mem_42 : _GEN_41; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_43 = 9'h2b == io_addra ? mem_43 : _GEN_42; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_44 = 9'h2c == io_addra ? mem_44 : _GEN_43; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_45 = 9'h2d == io_addra ? mem_45 : _GEN_44; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_46 = 9'h2e == io_addra ? mem_46 : _GEN_45; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_47 = 9'h2f == io_addra ? mem_47 : _GEN_46; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_48 = 9'h30 == io_addra ? mem_48 : _GEN_47; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_49 = 9'h31 == io_addra ? mem_49 : _GEN_48; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_50 = 9'h32 == io_addra ? mem_50 : _GEN_49; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_51 = 9'h33 == io_addra ? mem_51 : _GEN_50; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_52 = 9'h34 == io_addra ? mem_52 : _GEN_51; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_53 = 9'h35 == io_addra ? mem_53 : _GEN_52; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_54 = 9'h36 == io_addra ? mem_54 : _GEN_53; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_55 = 9'h37 == io_addra ? mem_55 : _GEN_54; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_56 = 9'h38 == io_addra ? mem_56 : _GEN_55; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_57 = 9'h39 == io_addra ? mem_57 : _GEN_56; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_58 = 9'h3a == io_addra ? mem_58 : _GEN_57; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_59 = 9'h3b == io_addra ? mem_59 : _GEN_58; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_60 = 9'h3c == io_addra ? mem_60 : _GEN_59; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_61 = 9'h3d == io_addra ? mem_61 : _GEN_60; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_62 = 9'h3e == io_addra ? mem_62 : _GEN_61; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_63 = 9'h3f == io_addra ? mem_63 : _GEN_62; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_64 = 9'h40 == io_addra ? mem_64 : _GEN_63; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_65 = 9'h41 == io_addra ? mem_65 : _GEN_64; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_66 = 9'h42 == io_addra ? mem_66 : _GEN_65; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_67 = 9'h43 == io_addra ? mem_67 : _GEN_66; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_68 = 9'h44 == io_addra ? mem_68 : _GEN_67; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_69 = 9'h45 == io_addra ? mem_69 : _GEN_68; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_70 = 9'h46 == io_addra ? mem_70 : _GEN_69; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_71 = 9'h47 == io_addra ? mem_71 : _GEN_70; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_72 = 9'h48 == io_addra ? mem_72 : _GEN_71; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_73 = 9'h49 == io_addra ? mem_73 : _GEN_72; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_74 = 9'h4a == io_addra ? mem_74 : _GEN_73; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_75 = 9'h4b == io_addra ? mem_75 : _GEN_74; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_76 = 9'h4c == io_addra ? mem_76 : _GEN_75; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_77 = 9'h4d == io_addra ? mem_77 : _GEN_76; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_78 = 9'h4e == io_addra ? mem_78 : _GEN_77; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_79 = 9'h4f == io_addra ? mem_79 : _GEN_78; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_80 = 9'h50 == io_addra ? mem_80 : _GEN_79; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_81 = 9'h51 == io_addra ? mem_81 : _GEN_80; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_82 = 9'h52 == io_addra ? mem_82 : _GEN_81; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_83 = 9'h53 == io_addra ? mem_83 : _GEN_82; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_84 = 9'h54 == io_addra ? mem_84 : _GEN_83; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_85 = 9'h55 == io_addra ? mem_85 : _GEN_84; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_86 = 9'h56 == io_addra ? mem_86 : _GEN_85; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_87 = 9'h57 == io_addra ? mem_87 : _GEN_86; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_88 = 9'h58 == io_addra ? mem_88 : _GEN_87; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_89 = 9'h59 == io_addra ? mem_89 : _GEN_88; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_90 = 9'h5a == io_addra ? mem_90 : _GEN_89; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_91 = 9'h5b == io_addra ? mem_91 : _GEN_90; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_92 = 9'h5c == io_addra ? mem_92 : _GEN_91; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_93 = 9'h5d == io_addra ? mem_93 : _GEN_92; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_94 = 9'h5e == io_addra ? mem_94 : _GEN_93; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_95 = 9'h5f == io_addra ? mem_95 : _GEN_94; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_96 = 9'h60 == io_addra ? mem_96 : _GEN_95; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_97 = 9'h61 == io_addra ? mem_97 : _GEN_96; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_98 = 9'h62 == io_addra ? mem_98 : _GEN_97; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_99 = 9'h63 == io_addra ? mem_99 : _GEN_98; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_100 = 9'h64 == io_addra ? mem_100 : _GEN_99; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_101 = 9'h65 == io_addra ? mem_101 : _GEN_100; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_102 = 9'h66 == io_addra ? mem_102 : _GEN_101; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_103 = 9'h67 == io_addra ? mem_103 : _GEN_102; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_104 = 9'h68 == io_addra ? mem_104 : _GEN_103; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_105 = 9'h69 == io_addra ? mem_105 : _GEN_104; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_106 = 9'h6a == io_addra ? mem_106 : _GEN_105; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_107 = 9'h6b == io_addra ? mem_107 : _GEN_106; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_108 = 9'h6c == io_addra ? mem_108 : _GEN_107; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_109 = 9'h6d == io_addra ? mem_109 : _GEN_108; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_110 = 9'h6e == io_addra ? mem_110 : _GEN_109; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_111 = 9'h6f == io_addra ? mem_111 : _GEN_110; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_112 = 9'h70 == io_addra ? mem_112 : _GEN_111; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_113 = 9'h71 == io_addra ? mem_113 : _GEN_112; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_114 = 9'h72 == io_addra ? mem_114 : _GEN_113; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_115 = 9'h73 == io_addra ? mem_115 : _GEN_114; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_116 = 9'h74 == io_addra ? mem_116 : _GEN_115; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_117 = 9'h75 == io_addra ? mem_117 : _GEN_116; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_118 = 9'h76 == io_addra ? mem_118 : _GEN_117; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_119 = 9'h77 == io_addra ? mem_119 : _GEN_118; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_120 = 9'h78 == io_addra ? mem_120 : _GEN_119; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_121 = 9'h79 == io_addra ? mem_121 : _GEN_120; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_122 = 9'h7a == io_addra ? mem_122 : _GEN_121; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_123 = 9'h7b == io_addra ? mem_123 : _GEN_122; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_124 = 9'h7c == io_addra ? mem_124 : _GEN_123; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_125 = 9'h7d == io_addra ? mem_125 : _GEN_124; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_126 = 9'h7e == io_addra ? mem_126 : _GEN_125; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_127 = 9'h7f == io_addra ? mem_127 : _GEN_126; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_128 = 9'h80 == io_addra ? mem_128 : _GEN_127; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_129 = 9'h81 == io_addra ? mem_129 : _GEN_128; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_130 = 9'h82 == io_addra ? mem_130 : _GEN_129; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_131 = 9'h83 == io_addra ? mem_131 : _GEN_130; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_132 = 9'h84 == io_addra ? mem_132 : _GEN_131; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_133 = 9'h85 == io_addra ? mem_133 : _GEN_132; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_134 = 9'h86 == io_addra ? mem_134 : _GEN_133; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_135 = 9'h87 == io_addra ? mem_135 : _GEN_134; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_136 = 9'h88 == io_addra ? mem_136 : _GEN_135; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_137 = 9'h89 == io_addra ? mem_137 : _GEN_136; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_138 = 9'h8a == io_addra ? mem_138 : _GEN_137; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_139 = 9'h8b == io_addra ? mem_139 : _GEN_138; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_140 = 9'h8c == io_addra ? mem_140 : _GEN_139; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_141 = 9'h8d == io_addra ? mem_141 : _GEN_140; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_142 = 9'h8e == io_addra ? mem_142 : _GEN_141; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_143 = 9'h8f == io_addra ? mem_143 : _GEN_142; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_144 = 9'h90 == io_addra ? mem_144 : _GEN_143; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_145 = 9'h91 == io_addra ? mem_145 : _GEN_144; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_146 = 9'h92 == io_addra ? mem_146 : _GEN_145; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_147 = 9'h93 == io_addra ? mem_147 : _GEN_146; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_148 = 9'h94 == io_addra ? mem_148 : _GEN_147; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_149 = 9'h95 == io_addra ? mem_149 : _GEN_148; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_150 = 9'h96 == io_addra ? mem_150 : _GEN_149; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_151 = 9'h97 == io_addra ? mem_151 : _GEN_150; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_152 = 9'h98 == io_addra ? mem_152 : _GEN_151; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_153 = 9'h99 == io_addra ? mem_153 : _GEN_152; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_154 = 9'h9a == io_addra ? mem_154 : _GEN_153; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_155 = 9'h9b == io_addra ? mem_155 : _GEN_154; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_156 = 9'h9c == io_addra ? mem_156 : _GEN_155; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_157 = 9'h9d == io_addra ? mem_157 : _GEN_156; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_158 = 9'h9e == io_addra ? mem_158 : _GEN_157; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_159 = 9'h9f == io_addra ? mem_159 : _GEN_158; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_160 = 9'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_161 = 9'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_162 = 9'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_163 = 9'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_164 = 9'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_165 = 9'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_166 = 9'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_167 = 9'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_168 = 9'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_169 = 9'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_170 = 9'haa == io_addra ? mem_170 : _GEN_169; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_171 = 9'hab == io_addra ? mem_171 : _GEN_170; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_172 = 9'hac == io_addra ? mem_172 : _GEN_171; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_173 = 9'had == io_addra ? mem_173 : _GEN_172; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_174 = 9'hae == io_addra ? mem_174 : _GEN_173; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_175 = 9'haf == io_addra ? mem_175 : _GEN_174; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_176 = 9'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_177 = 9'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_178 = 9'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_179 = 9'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_180 = 9'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_181 = 9'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_182 = 9'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_183 = 9'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_184 = 9'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_185 = 9'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_186 = 9'hba == io_addra ? mem_186 : _GEN_185; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_187 = 9'hbb == io_addra ? mem_187 : _GEN_186; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_188 = 9'hbc == io_addra ? mem_188 : _GEN_187; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_189 = 9'hbd == io_addra ? mem_189 : _GEN_188; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_190 = 9'hbe == io_addra ? mem_190 : _GEN_189; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_191 = 9'hbf == io_addra ? mem_191 : _GEN_190; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_192 = 9'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_193 = 9'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_194 = 9'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_195 = 9'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_196 = 9'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_197 = 9'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_198 = 9'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_199 = 9'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_200 = 9'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_201 = 9'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_202 = 9'hca == io_addra ? mem_202 : _GEN_201; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_203 = 9'hcb == io_addra ? mem_203 : _GEN_202; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_204 = 9'hcc == io_addra ? mem_204 : _GEN_203; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_205 = 9'hcd == io_addra ? mem_205 : _GEN_204; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_206 = 9'hce == io_addra ? mem_206 : _GEN_205; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_207 = 9'hcf == io_addra ? mem_207 : _GEN_206; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_208 = 9'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_209 = 9'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_210 = 9'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_211 = 9'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_212 = 9'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_213 = 9'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_214 = 9'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_215 = 9'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_216 = 9'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_217 = 9'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_218 = 9'hda == io_addra ? mem_218 : _GEN_217; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_219 = 9'hdb == io_addra ? mem_219 : _GEN_218; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_220 = 9'hdc == io_addra ? mem_220 : _GEN_219; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_221 = 9'hdd == io_addra ? mem_221 : _GEN_220; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_222 = 9'hde == io_addra ? mem_222 : _GEN_221; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_223 = 9'hdf == io_addra ? mem_223 : _GEN_222; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_224 = 9'he0 == io_addra ? mem_224 : _GEN_223; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_225 = 9'he1 == io_addra ? mem_225 : _GEN_224; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_226 = 9'he2 == io_addra ? mem_226 : _GEN_225; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_227 = 9'he3 == io_addra ? mem_227 : _GEN_226; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_228 = 9'he4 == io_addra ? mem_228 : _GEN_227; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_229 = 9'he5 == io_addra ? mem_229 : _GEN_228; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_230 = 9'he6 == io_addra ? mem_230 : _GEN_229; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_231 = 9'he7 == io_addra ? mem_231 : _GEN_230; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_232 = 9'he8 == io_addra ? mem_232 : _GEN_231; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_233 = 9'he9 == io_addra ? mem_233 : _GEN_232; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_234 = 9'hea == io_addra ? mem_234 : _GEN_233; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_235 = 9'heb == io_addra ? mem_235 : _GEN_234; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_236 = 9'hec == io_addra ? mem_236 : _GEN_235; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_237 = 9'hed == io_addra ? mem_237 : _GEN_236; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_238 = 9'hee == io_addra ? mem_238 : _GEN_237; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_239 = 9'hef == io_addra ? mem_239 : _GEN_238; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_240 = 9'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_241 = 9'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_242 = 9'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_243 = 9'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_244 = 9'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_245 = 9'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_246 = 9'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_247 = 9'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_248 = 9'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_249 = 9'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_250 = 9'hfa == io_addra ? mem_250 : _GEN_249; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_251 = 9'hfb == io_addra ? mem_251 : _GEN_250; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_252 = 9'hfc == io_addra ? mem_252 : _GEN_251; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_253 = 9'hfd == io_addra ? mem_253 : _GEN_252; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_254 = 9'hfe == io_addra ? mem_254 : _GEN_253; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_255 = 9'hff == io_addra ? mem_255 : _GEN_254; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_256 = 9'h100 == io_addra ? mem_256 : _GEN_255; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_257 = 9'h101 == io_addra ? mem_257 : _GEN_256; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_258 = 9'h102 == io_addra ? mem_258 : _GEN_257; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_259 = 9'h103 == io_addra ? mem_259 : _GEN_258; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_260 = 9'h104 == io_addra ? mem_260 : _GEN_259; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_261 = 9'h105 == io_addra ? mem_261 : _GEN_260; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_262 = 9'h106 == io_addra ? mem_262 : _GEN_261; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_263 = 9'h107 == io_addra ? mem_263 : _GEN_262; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_264 = 9'h108 == io_addra ? mem_264 : _GEN_263; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_265 = 9'h109 == io_addra ? mem_265 : _GEN_264; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_266 = 9'h10a == io_addra ? mem_266 : _GEN_265; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_267 = 9'h10b == io_addra ? mem_267 : _GEN_266; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_268 = 9'h10c == io_addra ? mem_268 : _GEN_267; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_269 = 9'h10d == io_addra ? mem_269 : _GEN_268; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_270 = 9'h10e == io_addra ? mem_270 : _GEN_269; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_271 = 9'h10f == io_addra ? mem_271 : _GEN_270; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_272 = 9'h110 == io_addra ? mem_272 : _GEN_271; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_273 = 9'h111 == io_addra ? mem_273 : _GEN_272; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_274 = 9'h112 == io_addra ? mem_274 : _GEN_273; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_275 = 9'h113 == io_addra ? mem_275 : _GEN_274; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_276 = 9'h114 == io_addra ? mem_276 : _GEN_275; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_277 = 9'h115 == io_addra ? mem_277 : _GEN_276; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_278 = 9'h116 == io_addra ? mem_278 : _GEN_277; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_279 = 9'h117 == io_addra ? mem_279 : _GEN_278; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_280 = 9'h118 == io_addra ? mem_280 : _GEN_279; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_281 = 9'h119 == io_addra ? mem_281 : _GEN_280; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_282 = 9'h11a == io_addra ? mem_282 : _GEN_281; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_283 = 9'h11b == io_addra ? mem_283 : _GEN_282; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_284 = 9'h11c == io_addra ? mem_284 : _GEN_283; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_285 = 9'h11d == io_addra ? mem_285 : _GEN_284; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_286 = 9'h11e == io_addra ? mem_286 : _GEN_285; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_287 = 9'h11f == io_addra ? mem_287 : _GEN_286; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_288 = 9'h120 == io_addra ? mem_288 : _GEN_287; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_289 = 9'h121 == io_addra ? mem_289 : _GEN_288; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_290 = 9'h122 == io_addra ? mem_290 : _GEN_289; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_291 = 9'h123 == io_addra ? mem_291 : _GEN_290; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_292 = 9'h124 == io_addra ? mem_292 : _GEN_291; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_293 = 9'h125 == io_addra ? mem_293 : _GEN_292; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_294 = 9'h126 == io_addra ? mem_294 : _GEN_293; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_295 = 9'h127 == io_addra ? mem_295 : _GEN_294; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_296 = 9'h128 == io_addra ? mem_296 : _GEN_295; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_297 = 9'h129 == io_addra ? mem_297 : _GEN_296; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_298 = 9'h12a == io_addra ? mem_298 : _GEN_297; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_299 = 9'h12b == io_addra ? mem_299 : _GEN_298; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_300 = 9'h12c == io_addra ? mem_300 : _GEN_299; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_301 = 9'h12d == io_addra ? mem_301 : _GEN_300; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_302 = 9'h12e == io_addra ? mem_302 : _GEN_301; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_303 = 9'h12f == io_addra ? mem_303 : _GEN_302; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_304 = 9'h130 == io_addra ? mem_304 : _GEN_303; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_305 = 9'h131 == io_addra ? mem_305 : _GEN_304; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_306 = 9'h132 == io_addra ? mem_306 : _GEN_305; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_307 = 9'h133 == io_addra ? mem_307 : _GEN_306; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_308 = 9'h134 == io_addra ? mem_308 : _GEN_307; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_309 = 9'h135 == io_addra ? mem_309 : _GEN_308; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_310 = 9'h136 == io_addra ? mem_310 : _GEN_309; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_311 = 9'h137 == io_addra ? mem_311 : _GEN_310; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_312 = 9'h138 == io_addra ? mem_312 : _GEN_311; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_313 = 9'h139 == io_addra ? mem_313 : _GEN_312; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_314 = 9'h13a == io_addra ? mem_314 : _GEN_313; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_315 = 9'h13b == io_addra ? mem_315 : _GEN_314; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_316 = 9'h13c == io_addra ? mem_316 : _GEN_315; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_317 = 9'h13d == io_addra ? mem_317 : _GEN_316; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_318 = 9'h13e == io_addra ? mem_318 : _GEN_317; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_319 = 9'h13f == io_addra ? mem_319 : _GEN_318; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_320 = 9'h140 == io_addra ? mem_320 : _GEN_319; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_321 = 9'h141 == io_addra ? mem_321 : _GEN_320; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_322 = 9'h142 == io_addra ? mem_322 : _GEN_321; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_323 = 9'h143 == io_addra ? mem_323 : _GEN_322; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_324 = 9'h144 == io_addra ? mem_324 : _GEN_323; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_325 = 9'h145 == io_addra ? mem_325 : _GEN_324; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_326 = 9'h146 == io_addra ? mem_326 : _GEN_325; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_327 = 9'h147 == io_addra ? mem_327 : _GEN_326; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_328 = 9'h148 == io_addra ? mem_328 : _GEN_327; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_329 = 9'h149 == io_addra ? mem_329 : _GEN_328; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_330 = 9'h14a == io_addra ? mem_330 : _GEN_329; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_331 = 9'h14b == io_addra ? mem_331 : _GEN_330; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_332 = 9'h14c == io_addra ? mem_332 : _GEN_331; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_333 = 9'h14d == io_addra ? mem_333 : _GEN_332; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_334 = 9'h14e == io_addra ? mem_334 : _GEN_333; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_335 = 9'h14f == io_addra ? mem_335 : _GEN_334; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_336 = 9'h150 == io_addra ? mem_336 : _GEN_335; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_337 = 9'h151 == io_addra ? mem_337 : _GEN_336; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_338 = 9'h152 == io_addra ? mem_338 : _GEN_337; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_339 = 9'h153 == io_addra ? mem_339 : _GEN_338; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_340 = 9'h154 == io_addra ? mem_340 : _GEN_339; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_341 = 9'h155 == io_addra ? mem_341 : _GEN_340; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_342 = 9'h156 == io_addra ? mem_342 : _GEN_341; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_343 = 9'h157 == io_addra ? mem_343 : _GEN_342; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_344 = 9'h158 == io_addra ? mem_344 : _GEN_343; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_345 = 9'h159 == io_addra ? mem_345 : _GEN_344; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_346 = 9'h15a == io_addra ? mem_346 : _GEN_345; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_347 = 9'h15b == io_addra ? mem_347 : _GEN_346; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_348 = 9'h15c == io_addra ? mem_348 : _GEN_347; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_349 = 9'h15d == io_addra ? mem_349 : _GEN_348; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_350 = 9'h15e == io_addra ? mem_350 : _GEN_349; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_351 = 9'h15f == io_addra ? mem_351 : _GEN_350; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_352 = 9'h160 == io_addra ? mem_352 : _GEN_351; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_353 = 9'h161 == io_addra ? mem_353 : _GEN_352; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_354 = 9'h162 == io_addra ? mem_354 : _GEN_353; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_355 = 9'h163 == io_addra ? mem_355 : _GEN_354; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_356 = 9'h164 == io_addra ? mem_356 : _GEN_355; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_357 = 9'h165 == io_addra ? mem_357 : _GEN_356; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_358 = 9'h166 == io_addra ? mem_358 : _GEN_357; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_359 = 9'h167 == io_addra ? mem_359 : _GEN_358; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_360 = 9'h168 == io_addra ? mem_360 : _GEN_359; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_361 = 9'h169 == io_addra ? mem_361 : _GEN_360; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_362 = 9'h16a == io_addra ? mem_362 : _GEN_361; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_363 = 9'h16b == io_addra ? mem_363 : _GEN_362; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_364 = 9'h16c == io_addra ? mem_364 : _GEN_363; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_365 = 9'h16d == io_addra ? mem_365 : _GEN_364; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_366 = 9'h16e == io_addra ? mem_366 : _GEN_365; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_367 = 9'h16f == io_addra ? mem_367 : _GEN_366; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_368 = 9'h170 == io_addra ? mem_368 : _GEN_367; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_369 = 9'h171 == io_addra ? mem_369 : _GEN_368; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_370 = 9'h172 == io_addra ? mem_370 : _GEN_369; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_371 = 9'h173 == io_addra ? mem_371 : _GEN_370; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_372 = 9'h174 == io_addra ? mem_372 : _GEN_371; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_373 = 9'h175 == io_addra ? mem_373 : _GEN_372; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_374 = 9'h176 == io_addra ? mem_374 : _GEN_373; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_375 = 9'h177 == io_addra ? mem_375 : _GEN_374; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_376 = 9'h178 == io_addra ? mem_376 : _GEN_375; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_377 = 9'h179 == io_addra ? mem_377 : _GEN_376; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_378 = 9'h17a == io_addra ? mem_378 : _GEN_377; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_379 = 9'h17b == io_addra ? mem_379 : _GEN_378; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_380 = 9'h17c == io_addra ? mem_380 : _GEN_379; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_381 = 9'h17d == io_addra ? mem_381 : _GEN_380; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_382 = 9'h17e == io_addra ? mem_382 : _GEN_381; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_383 = 9'h17f == io_addra ? mem_383 : _GEN_382; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_384 = 9'h180 == io_addra ? mem_384 : _GEN_383; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_385 = 9'h181 == io_addra ? mem_385 : _GEN_384; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_386 = 9'h182 == io_addra ? mem_386 : _GEN_385; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_387 = 9'h183 == io_addra ? mem_387 : _GEN_386; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_388 = 9'h184 == io_addra ? mem_388 : _GEN_387; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_389 = 9'h185 == io_addra ? mem_389 : _GEN_388; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_390 = 9'h186 == io_addra ? mem_390 : _GEN_389; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_391 = 9'h187 == io_addra ? mem_391 : _GEN_390; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_392 = 9'h188 == io_addra ? mem_392 : _GEN_391; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_393 = 9'h189 == io_addra ? mem_393 : _GEN_392; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_394 = 9'h18a == io_addra ? mem_394 : _GEN_393; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_395 = 9'h18b == io_addra ? mem_395 : _GEN_394; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_396 = 9'h18c == io_addra ? mem_396 : _GEN_395; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_397 = 9'h18d == io_addra ? mem_397 : _GEN_396; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_398 = 9'h18e == io_addra ? mem_398 : _GEN_397; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_399 = 9'h18f == io_addra ? mem_399 : _GEN_398; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_400 = 9'h190 == io_addra ? mem_400 : _GEN_399; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_401 = 9'h191 == io_addra ? mem_401 : _GEN_400; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_402 = 9'h192 == io_addra ? mem_402 : _GEN_401; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_403 = 9'h193 == io_addra ? mem_403 : _GEN_402; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_404 = 9'h194 == io_addra ? mem_404 : _GEN_403; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_405 = 9'h195 == io_addra ? mem_405 : _GEN_404; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_406 = 9'h196 == io_addra ? mem_406 : _GEN_405; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_407 = 9'h197 == io_addra ? mem_407 : _GEN_406; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_408 = 9'h198 == io_addra ? mem_408 : _GEN_407; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_409 = 9'h199 == io_addra ? mem_409 : _GEN_408; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_410 = 9'h19a == io_addra ? mem_410 : _GEN_409; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_411 = 9'h19b == io_addra ? mem_411 : _GEN_410; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_412 = 9'h19c == io_addra ? mem_412 : _GEN_411; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_413 = 9'h19d == io_addra ? mem_413 : _GEN_412; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_414 = 9'h19e == io_addra ? mem_414 : _GEN_413; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_415 = 9'h19f == io_addra ? mem_415 : _GEN_414; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_416 = 9'h1a0 == io_addra ? mem_416 : _GEN_415; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_417 = 9'h1a1 == io_addra ? mem_417 : _GEN_416; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_418 = 9'h1a2 == io_addra ? mem_418 : _GEN_417; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_419 = 9'h1a3 == io_addra ? mem_419 : _GEN_418; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_420 = 9'h1a4 == io_addra ? mem_420 : _GEN_419; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_421 = 9'h1a5 == io_addra ? mem_421 : _GEN_420; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_422 = 9'h1a6 == io_addra ? mem_422 : _GEN_421; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_423 = 9'h1a7 == io_addra ? mem_423 : _GEN_422; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_424 = 9'h1a8 == io_addra ? mem_424 : _GEN_423; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_425 = 9'h1a9 == io_addra ? mem_425 : _GEN_424; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_426 = 9'h1aa == io_addra ? mem_426 : _GEN_425; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_427 = 9'h1ab == io_addra ? mem_427 : _GEN_426; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_428 = 9'h1ac == io_addra ? mem_428 : _GEN_427; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_429 = 9'h1ad == io_addra ? mem_429 : _GEN_428; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_430 = 9'h1ae == io_addra ? mem_430 : _GEN_429; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_431 = 9'h1af == io_addra ? mem_431 : _GEN_430; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_432 = 9'h1b0 == io_addra ? mem_432 : _GEN_431; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_433 = 9'h1b1 == io_addra ? mem_433 : _GEN_432; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_434 = 9'h1b2 == io_addra ? mem_434 : _GEN_433; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_435 = 9'h1b3 == io_addra ? mem_435 : _GEN_434; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_436 = 9'h1b4 == io_addra ? mem_436 : _GEN_435; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_437 = 9'h1b5 == io_addra ? mem_437 : _GEN_436; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_438 = 9'h1b6 == io_addra ? mem_438 : _GEN_437; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_439 = 9'h1b7 == io_addra ? mem_439 : _GEN_438; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_440 = 9'h1b8 == io_addra ? mem_440 : _GEN_439; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_441 = 9'h1b9 == io_addra ? mem_441 : _GEN_440; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_442 = 9'h1ba == io_addra ? mem_442 : _GEN_441; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_443 = 9'h1bb == io_addra ? mem_443 : _GEN_442; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_444 = 9'h1bc == io_addra ? mem_444 : _GEN_443; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_445 = 9'h1bd == io_addra ? mem_445 : _GEN_444; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_446 = 9'h1be == io_addra ? mem_446 : _GEN_445; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_447 = 9'h1bf == io_addra ? mem_447 : _GEN_446; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_448 = 9'h1c0 == io_addra ? mem_448 : _GEN_447; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_449 = 9'h1c1 == io_addra ? mem_449 : _GEN_448; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_450 = 9'h1c2 == io_addra ? mem_450 : _GEN_449; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_451 = 9'h1c3 == io_addra ? mem_451 : _GEN_450; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_452 = 9'h1c4 == io_addra ? mem_452 : _GEN_451; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_453 = 9'h1c5 == io_addra ? mem_453 : _GEN_452; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_454 = 9'h1c6 == io_addra ? mem_454 : _GEN_453; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_455 = 9'h1c7 == io_addra ? mem_455 : _GEN_454; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_456 = 9'h1c8 == io_addra ? mem_456 : _GEN_455; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_457 = 9'h1c9 == io_addra ? mem_457 : _GEN_456; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_458 = 9'h1ca == io_addra ? mem_458 : _GEN_457; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_459 = 9'h1cb == io_addra ? mem_459 : _GEN_458; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_460 = 9'h1cc == io_addra ? mem_460 : _GEN_459; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_461 = 9'h1cd == io_addra ? mem_461 : _GEN_460; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_462 = 9'h1ce == io_addra ? mem_462 : _GEN_461; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_463 = 9'h1cf == io_addra ? mem_463 : _GEN_462; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_464 = 9'h1d0 == io_addra ? mem_464 : _GEN_463; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_465 = 9'h1d1 == io_addra ? mem_465 : _GEN_464; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_466 = 9'h1d2 == io_addra ? mem_466 : _GEN_465; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_467 = 9'h1d3 == io_addra ? mem_467 : _GEN_466; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_468 = 9'h1d4 == io_addra ? mem_468 : _GEN_467; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_469 = 9'h1d5 == io_addra ? mem_469 : _GEN_468; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_470 = 9'h1d6 == io_addra ? mem_470 : _GEN_469; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_471 = 9'h1d7 == io_addra ? mem_471 : _GEN_470; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_472 = 9'h1d8 == io_addra ? mem_472 : _GEN_471; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_473 = 9'h1d9 == io_addra ? mem_473 : _GEN_472; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_474 = 9'h1da == io_addra ? mem_474 : _GEN_473; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_475 = 9'h1db == io_addra ? mem_475 : _GEN_474; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_476 = 9'h1dc == io_addra ? mem_476 : _GEN_475; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_477 = 9'h1dd == io_addra ? mem_477 : _GEN_476; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_478 = 9'h1de == io_addra ? mem_478 : _GEN_477; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_479 = 9'h1df == io_addra ? mem_479 : _GEN_478; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_480 = 9'h1e0 == io_addra ? mem_480 : _GEN_479; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_481 = 9'h1e1 == io_addra ? mem_481 : _GEN_480; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_482 = 9'h1e2 == io_addra ? mem_482 : _GEN_481; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_483 = 9'h1e3 == io_addra ? mem_483 : _GEN_482; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_484 = 9'h1e4 == io_addra ? mem_484 : _GEN_483; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_485 = 9'h1e5 == io_addra ? mem_485 : _GEN_484; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_486 = 9'h1e6 == io_addra ? mem_486 : _GEN_485; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_487 = 9'h1e7 == io_addra ? mem_487 : _GEN_486; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_488 = 9'h1e8 == io_addra ? mem_488 : _GEN_487; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_489 = 9'h1e9 == io_addra ? mem_489 : _GEN_488; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_490 = 9'h1ea == io_addra ? mem_490 : _GEN_489; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_491 = 9'h1eb == io_addra ? mem_491 : _GEN_490; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_492 = 9'h1ec == io_addra ? mem_492 : _GEN_491; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_493 = 9'h1ed == io_addra ? mem_493 : _GEN_492; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_494 = 9'h1ee == io_addra ? mem_494 : _GEN_493; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_495 = 9'h1ef == io_addra ? mem_495 : _GEN_494; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_496 = 9'h1f0 == io_addra ? mem_496 : _GEN_495; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_497 = 9'h1f1 == io_addra ? mem_497 : _GEN_496; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_498 = 9'h1f2 == io_addra ? mem_498 : _GEN_497; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_499 = 9'h1f3 == io_addra ? mem_499 : _GEN_498; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_500 = 9'h1f4 == io_addra ? mem_500 : _GEN_499; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_501 = 9'h1f5 == io_addra ? mem_501 : _GEN_500; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_502 = 9'h1f6 == io_addra ? mem_502 : _GEN_501; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_503 = 9'h1f7 == io_addra ? mem_503 : _GEN_502; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_504 = 9'h1f8 == io_addra ? mem_504 : _GEN_503; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_505 = 9'h1f9 == io_addra ? mem_505 : _GEN_504; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_506 = 9'h1fa == io_addra ? mem_506 : _GEN_505; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [255:0] _GEN_507 = 9'h1fb == io_addra ? mem_507 : _GEN_506; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  assign io_douta = io_douta_REG; // @[RAMWrapper.scala 43:12]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_0 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_0 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_1 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_1 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_2 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_2 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_3 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_3 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_4 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_4 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_5 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_5 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_6 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_6 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_7 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_7 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_8 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_8 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_9 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_9 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_10 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_10 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_11 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_11 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_12 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_12 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_13 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_13 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_14 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_14 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_15 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_15 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_16 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_16 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_17 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_17 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_18 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_18 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_19 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_19 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_20 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_20 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_21 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_21 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_22 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_22 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_23 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_23 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_24 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_24 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_25 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_25 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_26 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_26 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_27 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_27 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_28 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_28 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_29 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_29 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_30 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_30 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_31 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_31 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_32 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h20 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_32 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_33 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h21 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_33 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_34 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h22 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_34 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_35 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h23 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_35 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_36 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h24 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_36 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_37 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h25 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_37 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_38 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h26 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_38 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_39 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h27 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_39 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_40 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h28 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_40 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_41 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h29 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_41 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_42 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_42 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_43 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_43 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_44 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_44 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_45 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_45 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_46 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_46 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_47 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_47 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_48 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h30 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_48 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_49 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h31 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_49 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_50 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h32 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_50 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_51 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h33 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_51 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_52 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h34 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_52 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_53 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h35 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_53 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_54 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h36 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_54 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_55 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h37 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_55 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_56 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h38 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_56 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_57 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h39 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_57 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_58 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_58 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_59 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_59 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_60 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_60 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_61 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_61 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_62 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_62 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_63 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_63 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_64 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h40 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_64 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_65 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h41 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_65 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_66 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h42 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_66 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_67 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h43 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_67 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_68 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h44 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_68 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_69 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h45 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_69 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_70 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h46 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_70 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_71 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h47 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_71 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_72 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h48 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_72 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_73 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h49 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_73 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_74 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_74 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_75 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_75 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_76 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_76 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_77 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_77 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_78 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_78 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_79 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_79 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_80 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h50 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_80 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_81 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h51 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_81 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_82 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h52 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_82 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_83 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h53 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_83 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_84 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h54 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_84 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_85 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h55 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_85 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_86 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h56 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_86 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_87 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h57 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_87 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_88 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h58 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_88 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_89 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h59 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_89 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_90 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_90 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_91 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_91 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_92 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_92 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_93 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_93 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_94 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_94 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_95 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_95 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_96 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h60 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_96 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_97 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h61 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_97 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_98 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h62 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_98 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_99 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h63 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_99 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_100 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h64 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_100 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_101 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h65 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_101 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_102 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h66 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_102 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_103 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h67 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_103 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_104 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h68 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_104 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_105 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h69 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_105 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_106 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_106 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_107 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_107 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_108 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_108 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_109 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_109 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_110 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_110 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_111 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_111 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_112 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h70 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_112 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_113 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h71 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_113 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_114 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h72 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_114 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_115 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h73 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_115 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_116 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h74 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_116 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_117 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h75 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_117 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_118 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h76 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_118 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_119 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h77 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_119 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_120 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h78 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_120 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_121 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h79 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_121 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_122 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_122 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_123 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_123 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_124 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_124 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_125 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_125 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_126 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_126 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_127 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_127 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_128 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h80 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_128 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_129 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h81 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_129 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_130 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h82 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_130 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_131 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h83 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_131 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_132 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h84 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_132 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_133 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h85 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_133 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_134 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h86 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_134 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_135 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h87 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_135 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_136 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h88 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_136 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_137 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h89 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_137 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_138 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_138 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_139 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_139 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_140 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_140 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_141 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_141 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_142 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_142 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_143 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_143 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_144 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h90 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_144 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_145 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h91 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_145 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_146 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h92 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_146 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_147 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h93 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_147 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_148 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h94 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_148 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_149 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h95 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_149 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_150 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h96 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_150 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_151 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h97 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_151 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_152 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h98 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_152 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_153 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h99 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_153 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_154 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_154 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_155 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_155 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_156 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_156 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_157 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_157 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_158 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_158 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_159 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_159 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_160 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_160 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_161 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_161 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_162 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_162 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_163 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_163 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_164 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_164 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_165 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_165 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_166 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_166 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_167 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_167 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_168 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_168 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_169 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_169 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_170 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'haa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_170 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_171 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hab == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_171 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_172 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hac == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_172 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_173 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'had == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_173 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_174 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hae == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_174 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_175 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'haf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_175 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_176 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_176 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_177 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_177 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_178 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_178 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_179 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_179 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_180 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_180 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_181 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_181 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_182 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_182 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_183 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_183 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_184 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_184 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_185 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_185 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_186 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hba == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_186 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_187 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_187 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_188 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_188 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_189 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_189 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_190 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_190 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_191 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_191 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_192 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_192 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_193 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_193 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_194 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_194 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_195 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_195 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_196 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_196 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_197 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_197 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_198 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_198 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_199 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_199 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_200 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_200 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_201 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_201 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_202 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hca == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_202 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_203 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_203 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_204 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_204 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_205 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_205 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_206 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hce == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_206 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_207 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_207 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_208 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_208 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_209 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_209 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_210 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_210 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_211 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_211 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_212 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_212 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_213 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_213 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_214 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_214 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_215 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_215 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_216 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_216 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_217 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_217 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_218 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hda == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_218 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_219 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_219 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_220 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_220 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_221 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_221 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_222 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hde == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_222 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_223 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_223 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_224 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_224 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_225 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_225 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_226 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_226 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_227 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_227 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_228 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_228 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_229 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_229 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_230 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_230 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_231 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_231 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_232 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_232 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_233 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_233 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_234 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hea == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_234 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_235 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'heb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_235 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_236 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hec == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_236 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_237 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hed == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_237 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_238 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hee == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_238 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_239 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hef == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_239 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_240 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_240 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_241 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_241 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_242 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_242 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_243 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_243 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_244 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_244 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_245 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_245 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_246 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_246 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_247 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_247 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_248 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_248 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_249 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_249 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_250 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_250 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_251 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_251 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_252 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_252 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_253 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_253 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_254 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_254 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_255 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hff == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_255 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_256 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h100 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_256 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_257 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h101 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_257 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_258 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h102 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_258 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_259 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h103 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_259 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_260 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h104 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_260 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_261 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h105 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_261 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_262 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h106 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_262 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_263 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h107 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_263 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_264 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h108 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_264 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_265 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h109 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_265 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_266 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_266 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_267 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_267 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_268 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_268 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_269 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_269 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_270 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_270 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_271 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_271 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_272 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h110 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_272 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_273 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h111 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_273 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_274 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h112 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_274 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_275 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h113 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_275 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_276 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h114 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_276 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_277 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h115 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_277 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_278 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h116 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_278 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_279 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h117 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_279 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_280 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h118 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_280 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_281 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h119 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_281 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_282 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_282 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_283 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_283 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_284 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_284 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_285 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_285 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_286 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_286 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_287 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_287 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_288 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h120 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_288 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_289 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h121 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_289 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_290 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h122 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_290 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_291 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h123 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_291 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_292 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h124 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_292 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_293 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h125 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_293 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_294 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h126 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_294 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_295 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h127 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_295 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_296 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h128 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_296 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_297 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h129 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_297 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_298 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_298 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_299 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_299 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_300 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_300 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_301 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_301 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_302 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_302 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_303 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_303 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_304 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h130 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_304 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_305 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h131 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_305 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_306 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h132 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_306 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_307 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h133 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_307 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_308 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h134 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_308 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_309 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h135 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_309 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_310 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h136 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_310 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_311 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h137 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_311 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_312 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h138 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_312 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_313 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h139 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_313 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_314 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_314 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_315 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_315 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_316 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_316 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_317 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_317 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_318 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_318 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_319 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_319 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_320 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h140 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_320 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_321 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h141 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_321 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_322 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h142 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_322 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_323 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h143 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_323 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_324 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h144 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_324 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_325 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h145 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_325 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_326 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h146 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_326 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_327 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h147 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_327 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_328 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h148 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_328 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_329 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h149 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_329 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_330 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_330 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_331 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_331 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_332 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_332 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_333 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_333 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_334 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_334 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_335 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_335 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_336 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h150 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_336 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_337 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h151 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_337 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_338 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h152 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_338 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_339 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h153 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_339 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_340 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h154 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_340 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_341 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h155 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_341 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_342 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h156 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_342 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_343 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h157 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_343 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_344 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h158 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_344 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_345 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h159 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_345 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_346 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_346 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_347 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_347 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_348 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_348 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_349 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_349 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_350 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_350 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_351 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_351 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_352 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h160 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_352 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_353 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h161 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_353 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_354 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h162 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_354 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_355 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h163 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_355 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_356 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h164 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_356 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_357 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h165 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_357 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_358 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h166 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_358 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_359 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h167 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_359 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_360 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h168 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_360 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_361 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h169 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_361 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_362 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_362 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_363 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_363 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_364 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_364 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_365 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_365 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_366 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_366 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_367 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_367 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_368 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h170 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_368 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_369 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h171 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_369 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_370 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h172 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_370 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_371 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h173 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_371 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_372 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h174 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_372 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_373 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h175 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_373 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_374 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h176 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_374 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_375 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h177 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_375 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_376 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h178 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_376 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_377 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h179 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_377 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_378 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_378 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_379 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_379 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_380 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_380 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_381 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_381 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_382 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_382 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_383 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_383 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_384 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h180 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_384 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_385 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h181 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_385 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_386 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h182 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_386 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_387 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h183 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_387 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_388 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h184 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_388 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_389 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h185 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_389 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_390 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h186 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_390 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_391 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h187 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_391 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_392 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h188 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_392 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_393 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h189 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_393 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_394 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_394 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_395 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_395 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_396 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_396 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_397 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_397 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_398 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_398 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_399 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_399 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_400 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h190 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_400 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_401 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h191 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_401 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_402 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h192 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_402 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_403 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h193 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_403 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_404 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h194 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_404 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_405 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h195 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_405 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_406 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h196 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_406 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_407 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h197 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_407 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_408 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h198 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_408 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_409 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h199 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_409 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_410 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_410 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_411 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_411 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_412 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_412 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_413 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_413 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_414 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_414 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_415 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_415 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_416 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_416 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_417 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_417 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_418 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_418 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_419 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_419 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_420 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_420 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_421 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_421 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_422 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_422 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_423 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_423 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_424 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_424 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_425 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_425 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_426 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1aa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_426 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_427 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ab == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_427 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_428 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ac == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_428 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_429 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ad == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_429 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_430 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ae == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_430 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_431 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1af == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_431 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_432 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_432 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_433 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_433 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_434 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_434 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_435 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_435 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_436 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_436 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_437 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_437 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_438 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_438 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_439 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_439 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_440 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_440 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_441 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_441 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_442 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ba == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_442 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_443 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_443 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_444 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_444 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_445 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_445 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_446 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1be == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_446 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_447 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_447 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_448 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_448 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_449 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_449 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_450 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_450 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_451 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_451 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_452 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_452 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_453 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_453 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_454 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_454 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_455 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_455 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_456 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_456 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_457 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_457 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_458 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ca == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_458 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_459 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_459 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_460 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_460 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_461 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_461 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_462 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ce == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_462 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_463 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_463 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_464 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_464 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_465 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_465 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_466 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_466 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_467 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_467 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_468 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_468 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_469 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_469 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_470 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_470 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_471 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_471 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_472 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_472 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_473 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_473 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_474 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1da == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_474 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_475 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1db == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_475 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_476 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1dc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_476 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_477 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1dd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_477 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_478 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1de == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_478 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_479 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1df == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_479 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_480 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_480 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_481 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_481 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_482 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_482 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_483 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_483 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_484 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_484 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_485 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_485 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_486 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_486 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_487 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_487 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_488 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_488 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_489 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_489 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_490 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ea == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_490 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_491 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1eb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_491 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_492 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ec == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_492 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_493 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ed == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_493 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_494 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ee == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_494 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_495 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ef == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_495 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_496 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_496 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_497 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_497 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_498 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_498 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_499 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_499 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_500 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_500 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_501 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_501 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_502 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_502 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_503 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_503 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_504 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_504 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_505 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_505 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_506 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_506 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_507 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_507 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_508 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_508 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_509 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_509 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_510 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_510 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_511 <= 256'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ff == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_511 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (9'h1ff == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_511; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fe == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_510; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fd == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_509; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fc == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_508; // @[RAMWrapper.scala 43:22]
    end else begin
      io_douta_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  mem_0 = _RAND_0[255:0];
  _RAND_1 = {8{`RANDOM}};
  mem_1 = _RAND_1[255:0];
  _RAND_2 = {8{`RANDOM}};
  mem_2 = _RAND_2[255:0];
  _RAND_3 = {8{`RANDOM}};
  mem_3 = _RAND_3[255:0];
  _RAND_4 = {8{`RANDOM}};
  mem_4 = _RAND_4[255:0];
  _RAND_5 = {8{`RANDOM}};
  mem_5 = _RAND_5[255:0];
  _RAND_6 = {8{`RANDOM}};
  mem_6 = _RAND_6[255:0];
  _RAND_7 = {8{`RANDOM}};
  mem_7 = _RAND_7[255:0];
  _RAND_8 = {8{`RANDOM}};
  mem_8 = _RAND_8[255:0];
  _RAND_9 = {8{`RANDOM}};
  mem_9 = _RAND_9[255:0];
  _RAND_10 = {8{`RANDOM}};
  mem_10 = _RAND_10[255:0];
  _RAND_11 = {8{`RANDOM}};
  mem_11 = _RAND_11[255:0];
  _RAND_12 = {8{`RANDOM}};
  mem_12 = _RAND_12[255:0];
  _RAND_13 = {8{`RANDOM}};
  mem_13 = _RAND_13[255:0];
  _RAND_14 = {8{`RANDOM}};
  mem_14 = _RAND_14[255:0];
  _RAND_15 = {8{`RANDOM}};
  mem_15 = _RAND_15[255:0];
  _RAND_16 = {8{`RANDOM}};
  mem_16 = _RAND_16[255:0];
  _RAND_17 = {8{`RANDOM}};
  mem_17 = _RAND_17[255:0];
  _RAND_18 = {8{`RANDOM}};
  mem_18 = _RAND_18[255:0];
  _RAND_19 = {8{`RANDOM}};
  mem_19 = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  mem_20 = _RAND_20[255:0];
  _RAND_21 = {8{`RANDOM}};
  mem_21 = _RAND_21[255:0];
  _RAND_22 = {8{`RANDOM}};
  mem_22 = _RAND_22[255:0];
  _RAND_23 = {8{`RANDOM}};
  mem_23 = _RAND_23[255:0];
  _RAND_24 = {8{`RANDOM}};
  mem_24 = _RAND_24[255:0];
  _RAND_25 = {8{`RANDOM}};
  mem_25 = _RAND_25[255:0];
  _RAND_26 = {8{`RANDOM}};
  mem_26 = _RAND_26[255:0];
  _RAND_27 = {8{`RANDOM}};
  mem_27 = _RAND_27[255:0];
  _RAND_28 = {8{`RANDOM}};
  mem_28 = _RAND_28[255:0];
  _RAND_29 = {8{`RANDOM}};
  mem_29 = _RAND_29[255:0];
  _RAND_30 = {8{`RANDOM}};
  mem_30 = _RAND_30[255:0];
  _RAND_31 = {8{`RANDOM}};
  mem_31 = _RAND_31[255:0];
  _RAND_32 = {8{`RANDOM}};
  mem_32 = _RAND_32[255:0];
  _RAND_33 = {8{`RANDOM}};
  mem_33 = _RAND_33[255:0];
  _RAND_34 = {8{`RANDOM}};
  mem_34 = _RAND_34[255:0];
  _RAND_35 = {8{`RANDOM}};
  mem_35 = _RAND_35[255:0];
  _RAND_36 = {8{`RANDOM}};
  mem_36 = _RAND_36[255:0];
  _RAND_37 = {8{`RANDOM}};
  mem_37 = _RAND_37[255:0];
  _RAND_38 = {8{`RANDOM}};
  mem_38 = _RAND_38[255:0];
  _RAND_39 = {8{`RANDOM}};
  mem_39 = _RAND_39[255:0];
  _RAND_40 = {8{`RANDOM}};
  mem_40 = _RAND_40[255:0];
  _RAND_41 = {8{`RANDOM}};
  mem_41 = _RAND_41[255:0];
  _RAND_42 = {8{`RANDOM}};
  mem_42 = _RAND_42[255:0];
  _RAND_43 = {8{`RANDOM}};
  mem_43 = _RAND_43[255:0];
  _RAND_44 = {8{`RANDOM}};
  mem_44 = _RAND_44[255:0];
  _RAND_45 = {8{`RANDOM}};
  mem_45 = _RAND_45[255:0];
  _RAND_46 = {8{`RANDOM}};
  mem_46 = _RAND_46[255:0];
  _RAND_47 = {8{`RANDOM}};
  mem_47 = _RAND_47[255:0];
  _RAND_48 = {8{`RANDOM}};
  mem_48 = _RAND_48[255:0];
  _RAND_49 = {8{`RANDOM}};
  mem_49 = _RAND_49[255:0];
  _RAND_50 = {8{`RANDOM}};
  mem_50 = _RAND_50[255:0];
  _RAND_51 = {8{`RANDOM}};
  mem_51 = _RAND_51[255:0];
  _RAND_52 = {8{`RANDOM}};
  mem_52 = _RAND_52[255:0];
  _RAND_53 = {8{`RANDOM}};
  mem_53 = _RAND_53[255:0];
  _RAND_54 = {8{`RANDOM}};
  mem_54 = _RAND_54[255:0];
  _RAND_55 = {8{`RANDOM}};
  mem_55 = _RAND_55[255:0];
  _RAND_56 = {8{`RANDOM}};
  mem_56 = _RAND_56[255:0];
  _RAND_57 = {8{`RANDOM}};
  mem_57 = _RAND_57[255:0];
  _RAND_58 = {8{`RANDOM}};
  mem_58 = _RAND_58[255:0];
  _RAND_59 = {8{`RANDOM}};
  mem_59 = _RAND_59[255:0];
  _RAND_60 = {8{`RANDOM}};
  mem_60 = _RAND_60[255:0];
  _RAND_61 = {8{`RANDOM}};
  mem_61 = _RAND_61[255:0];
  _RAND_62 = {8{`RANDOM}};
  mem_62 = _RAND_62[255:0];
  _RAND_63 = {8{`RANDOM}};
  mem_63 = _RAND_63[255:0];
  _RAND_64 = {8{`RANDOM}};
  mem_64 = _RAND_64[255:0];
  _RAND_65 = {8{`RANDOM}};
  mem_65 = _RAND_65[255:0];
  _RAND_66 = {8{`RANDOM}};
  mem_66 = _RAND_66[255:0];
  _RAND_67 = {8{`RANDOM}};
  mem_67 = _RAND_67[255:0];
  _RAND_68 = {8{`RANDOM}};
  mem_68 = _RAND_68[255:0];
  _RAND_69 = {8{`RANDOM}};
  mem_69 = _RAND_69[255:0];
  _RAND_70 = {8{`RANDOM}};
  mem_70 = _RAND_70[255:0];
  _RAND_71 = {8{`RANDOM}};
  mem_71 = _RAND_71[255:0];
  _RAND_72 = {8{`RANDOM}};
  mem_72 = _RAND_72[255:0];
  _RAND_73 = {8{`RANDOM}};
  mem_73 = _RAND_73[255:0];
  _RAND_74 = {8{`RANDOM}};
  mem_74 = _RAND_74[255:0];
  _RAND_75 = {8{`RANDOM}};
  mem_75 = _RAND_75[255:0];
  _RAND_76 = {8{`RANDOM}};
  mem_76 = _RAND_76[255:0];
  _RAND_77 = {8{`RANDOM}};
  mem_77 = _RAND_77[255:0];
  _RAND_78 = {8{`RANDOM}};
  mem_78 = _RAND_78[255:0];
  _RAND_79 = {8{`RANDOM}};
  mem_79 = _RAND_79[255:0];
  _RAND_80 = {8{`RANDOM}};
  mem_80 = _RAND_80[255:0];
  _RAND_81 = {8{`RANDOM}};
  mem_81 = _RAND_81[255:0];
  _RAND_82 = {8{`RANDOM}};
  mem_82 = _RAND_82[255:0];
  _RAND_83 = {8{`RANDOM}};
  mem_83 = _RAND_83[255:0];
  _RAND_84 = {8{`RANDOM}};
  mem_84 = _RAND_84[255:0];
  _RAND_85 = {8{`RANDOM}};
  mem_85 = _RAND_85[255:0];
  _RAND_86 = {8{`RANDOM}};
  mem_86 = _RAND_86[255:0];
  _RAND_87 = {8{`RANDOM}};
  mem_87 = _RAND_87[255:0];
  _RAND_88 = {8{`RANDOM}};
  mem_88 = _RAND_88[255:0];
  _RAND_89 = {8{`RANDOM}};
  mem_89 = _RAND_89[255:0];
  _RAND_90 = {8{`RANDOM}};
  mem_90 = _RAND_90[255:0];
  _RAND_91 = {8{`RANDOM}};
  mem_91 = _RAND_91[255:0];
  _RAND_92 = {8{`RANDOM}};
  mem_92 = _RAND_92[255:0];
  _RAND_93 = {8{`RANDOM}};
  mem_93 = _RAND_93[255:0];
  _RAND_94 = {8{`RANDOM}};
  mem_94 = _RAND_94[255:0];
  _RAND_95 = {8{`RANDOM}};
  mem_95 = _RAND_95[255:0];
  _RAND_96 = {8{`RANDOM}};
  mem_96 = _RAND_96[255:0];
  _RAND_97 = {8{`RANDOM}};
  mem_97 = _RAND_97[255:0];
  _RAND_98 = {8{`RANDOM}};
  mem_98 = _RAND_98[255:0];
  _RAND_99 = {8{`RANDOM}};
  mem_99 = _RAND_99[255:0];
  _RAND_100 = {8{`RANDOM}};
  mem_100 = _RAND_100[255:0];
  _RAND_101 = {8{`RANDOM}};
  mem_101 = _RAND_101[255:0];
  _RAND_102 = {8{`RANDOM}};
  mem_102 = _RAND_102[255:0];
  _RAND_103 = {8{`RANDOM}};
  mem_103 = _RAND_103[255:0];
  _RAND_104 = {8{`RANDOM}};
  mem_104 = _RAND_104[255:0];
  _RAND_105 = {8{`RANDOM}};
  mem_105 = _RAND_105[255:0];
  _RAND_106 = {8{`RANDOM}};
  mem_106 = _RAND_106[255:0];
  _RAND_107 = {8{`RANDOM}};
  mem_107 = _RAND_107[255:0];
  _RAND_108 = {8{`RANDOM}};
  mem_108 = _RAND_108[255:0];
  _RAND_109 = {8{`RANDOM}};
  mem_109 = _RAND_109[255:0];
  _RAND_110 = {8{`RANDOM}};
  mem_110 = _RAND_110[255:0];
  _RAND_111 = {8{`RANDOM}};
  mem_111 = _RAND_111[255:0];
  _RAND_112 = {8{`RANDOM}};
  mem_112 = _RAND_112[255:0];
  _RAND_113 = {8{`RANDOM}};
  mem_113 = _RAND_113[255:0];
  _RAND_114 = {8{`RANDOM}};
  mem_114 = _RAND_114[255:0];
  _RAND_115 = {8{`RANDOM}};
  mem_115 = _RAND_115[255:0];
  _RAND_116 = {8{`RANDOM}};
  mem_116 = _RAND_116[255:0];
  _RAND_117 = {8{`RANDOM}};
  mem_117 = _RAND_117[255:0];
  _RAND_118 = {8{`RANDOM}};
  mem_118 = _RAND_118[255:0];
  _RAND_119 = {8{`RANDOM}};
  mem_119 = _RAND_119[255:0];
  _RAND_120 = {8{`RANDOM}};
  mem_120 = _RAND_120[255:0];
  _RAND_121 = {8{`RANDOM}};
  mem_121 = _RAND_121[255:0];
  _RAND_122 = {8{`RANDOM}};
  mem_122 = _RAND_122[255:0];
  _RAND_123 = {8{`RANDOM}};
  mem_123 = _RAND_123[255:0];
  _RAND_124 = {8{`RANDOM}};
  mem_124 = _RAND_124[255:0];
  _RAND_125 = {8{`RANDOM}};
  mem_125 = _RAND_125[255:0];
  _RAND_126 = {8{`RANDOM}};
  mem_126 = _RAND_126[255:0];
  _RAND_127 = {8{`RANDOM}};
  mem_127 = _RAND_127[255:0];
  _RAND_128 = {8{`RANDOM}};
  mem_128 = _RAND_128[255:0];
  _RAND_129 = {8{`RANDOM}};
  mem_129 = _RAND_129[255:0];
  _RAND_130 = {8{`RANDOM}};
  mem_130 = _RAND_130[255:0];
  _RAND_131 = {8{`RANDOM}};
  mem_131 = _RAND_131[255:0];
  _RAND_132 = {8{`RANDOM}};
  mem_132 = _RAND_132[255:0];
  _RAND_133 = {8{`RANDOM}};
  mem_133 = _RAND_133[255:0];
  _RAND_134 = {8{`RANDOM}};
  mem_134 = _RAND_134[255:0];
  _RAND_135 = {8{`RANDOM}};
  mem_135 = _RAND_135[255:0];
  _RAND_136 = {8{`RANDOM}};
  mem_136 = _RAND_136[255:0];
  _RAND_137 = {8{`RANDOM}};
  mem_137 = _RAND_137[255:0];
  _RAND_138 = {8{`RANDOM}};
  mem_138 = _RAND_138[255:0];
  _RAND_139 = {8{`RANDOM}};
  mem_139 = _RAND_139[255:0];
  _RAND_140 = {8{`RANDOM}};
  mem_140 = _RAND_140[255:0];
  _RAND_141 = {8{`RANDOM}};
  mem_141 = _RAND_141[255:0];
  _RAND_142 = {8{`RANDOM}};
  mem_142 = _RAND_142[255:0];
  _RAND_143 = {8{`RANDOM}};
  mem_143 = _RAND_143[255:0];
  _RAND_144 = {8{`RANDOM}};
  mem_144 = _RAND_144[255:0];
  _RAND_145 = {8{`RANDOM}};
  mem_145 = _RAND_145[255:0];
  _RAND_146 = {8{`RANDOM}};
  mem_146 = _RAND_146[255:0];
  _RAND_147 = {8{`RANDOM}};
  mem_147 = _RAND_147[255:0];
  _RAND_148 = {8{`RANDOM}};
  mem_148 = _RAND_148[255:0];
  _RAND_149 = {8{`RANDOM}};
  mem_149 = _RAND_149[255:0];
  _RAND_150 = {8{`RANDOM}};
  mem_150 = _RAND_150[255:0];
  _RAND_151 = {8{`RANDOM}};
  mem_151 = _RAND_151[255:0];
  _RAND_152 = {8{`RANDOM}};
  mem_152 = _RAND_152[255:0];
  _RAND_153 = {8{`RANDOM}};
  mem_153 = _RAND_153[255:0];
  _RAND_154 = {8{`RANDOM}};
  mem_154 = _RAND_154[255:0];
  _RAND_155 = {8{`RANDOM}};
  mem_155 = _RAND_155[255:0];
  _RAND_156 = {8{`RANDOM}};
  mem_156 = _RAND_156[255:0];
  _RAND_157 = {8{`RANDOM}};
  mem_157 = _RAND_157[255:0];
  _RAND_158 = {8{`RANDOM}};
  mem_158 = _RAND_158[255:0];
  _RAND_159 = {8{`RANDOM}};
  mem_159 = _RAND_159[255:0];
  _RAND_160 = {8{`RANDOM}};
  mem_160 = _RAND_160[255:0];
  _RAND_161 = {8{`RANDOM}};
  mem_161 = _RAND_161[255:0];
  _RAND_162 = {8{`RANDOM}};
  mem_162 = _RAND_162[255:0];
  _RAND_163 = {8{`RANDOM}};
  mem_163 = _RAND_163[255:0];
  _RAND_164 = {8{`RANDOM}};
  mem_164 = _RAND_164[255:0];
  _RAND_165 = {8{`RANDOM}};
  mem_165 = _RAND_165[255:0];
  _RAND_166 = {8{`RANDOM}};
  mem_166 = _RAND_166[255:0];
  _RAND_167 = {8{`RANDOM}};
  mem_167 = _RAND_167[255:0];
  _RAND_168 = {8{`RANDOM}};
  mem_168 = _RAND_168[255:0];
  _RAND_169 = {8{`RANDOM}};
  mem_169 = _RAND_169[255:0];
  _RAND_170 = {8{`RANDOM}};
  mem_170 = _RAND_170[255:0];
  _RAND_171 = {8{`RANDOM}};
  mem_171 = _RAND_171[255:0];
  _RAND_172 = {8{`RANDOM}};
  mem_172 = _RAND_172[255:0];
  _RAND_173 = {8{`RANDOM}};
  mem_173 = _RAND_173[255:0];
  _RAND_174 = {8{`RANDOM}};
  mem_174 = _RAND_174[255:0];
  _RAND_175 = {8{`RANDOM}};
  mem_175 = _RAND_175[255:0];
  _RAND_176 = {8{`RANDOM}};
  mem_176 = _RAND_176[255:0];
  _RAND_177 = {8{`RANDOM}};
  mem_177 = _RAND_177[255:0];
  _RAND_178 = {8{`RANDOM}};
  mem_178 = _RAND_178[255:0];
  _RAND_179 = {8{`RANDOM}};
  mem_179 = _RAND_179[255:0];
  _RAND_180 = {8{`RANDOM}};
  mem_180 = _RAND_180[255:0];
  _RAND_181 = {8{`RANDOM}};
  mem_181 = _RAND_181[255:0];
  _RAND_182 = {8{`RANDOM}};
  mem_182 = _RAND_182[255:0];
  _RAND_183 = {8{`RANDOM}};
  mem_183 = _RAND_183[255:0];
  _RAND_184 = {8{`RANDOM}};
  mem_184 = _RAND_184[255:0];
  _RAND_185 = {8{`RANDOM}};
  mem_185 = _RAND_185[255:0];
  _RAND_186 = {8{`RANDOM}};
  mem_186 = _RAND_186[255:0];
  _RAND_187 = {8{`RANDOM}};
  mem_187 = _RAND_187[255:0];
  _RAND_188 = {8{`RANDOM}};
  mem_188 = _RAND_188[255:0];
  _RAND_189 = {8{`RANDOM}};
  mem_189 = _RAND_189[255:0];
  _RAND_190 = {8{`RANDOM}};
  mem_190 = _RAND_190[255:0];
  _RAND_191 = {8{`RANDOM}};
  mem_191 = _RAND_191[255:0];
  _RAND_192 = {8{`RANDOM}};
  mem_192 = _RAND_192[255:0];
  _RAND_193 = {8{`RANDOM}};
  mem_193 = _RAND_193[255:0];
  _RAND_194 = {8{`RANDOM}};
  mem_194 = _RAND_194[255:0];
  _RAND_195 = {8{`RANDOM}};
  mem_195 = _RAND_195[255:0];
  _RAND_196 = {8{`RANDOM}};
  mem_196 = _RAND_196[255:0];
  _RAND_197 = {8{`RANDOM}};
  mem_197 = _RAND_197[255:0];
  _RAND_198 = {8{`RANDOM}};
  mem_198 = _RAND_198[255:0];
  _RAND_199 = {8{`RANDOM}};
  mem_199 = _RAND_199[255:0];
  _RAND_200 = {8{`RANDOM}};
  mem_200 = _RAND_200[255:0];
  _RAND_201 = {8{`RANDOM}};
  mem_201 = _RAND_201[255:0];
  _RAND_202 = {8{`RANDOM}};
  mem_202 = _RAND_202[255:0];
  _RAND_203 = {8{`RANDOM}};
  mem_203 = _RAND_203[255:0];
  _RAND_204 = {8{`RANDOM}};
  mem_204 = _RAND_204[255:0];
  _RAND_205 = {8{`RANDOM}};
  mem_205 = _RAND_205[255:0];
  _RAND_206 = {8{`RANDOM}};
  mem_206 = _RAND_206[255:0];
  _RAND_207 = {8{`RANDOM}};
  mem_207 = _RAND_207[255:0];
  _RAND_208 = {8{`RANDOM}};
  mem_208 = _RAND_208[255:0];
  _RAND_209 = {8{`RANDOM}};
  mem_209 = _RAND_209[255:0];
  _RAND_210 = {8{`RANDOM}};
  mem_210 = _RAND_210[255:0];
  _RAND_211 = {8{`RANDOM}};
  mem_211 = _RAND_211[255:0];
  _RAND_212 = {8{`RANDOM}};
  mem_212 = _RAND_212[255:0];
  _RAND_213 = {8{`RANDOM}};
  mem_213 = _RAND_213[255:0];
  _RAND_214 = {8{`RANDOM}};
  mem_214 = _RAND_214[255:0];
  _RAND_215 = {8{`RANDOM}};
  mem_215 = _RAND_215[255:0];
  _RAND_216 = {8{`RANDOM}};
  mem_216 = _RAND_216[255:0];
  _RAND_217 = {8{`RANDOM}};
  mem_217 = _RAND_217[255:0];
  _RAND_218 = {8{`RANDOM}};
  mem_218 = _RAND_218[255:0];
  _RAND_219 = {8{`RANDOM}};
  mem_219 = _RAND_219[255:0];
  _RAND_220 = {8{`RANDOM}};
  mem_220 = _RAND_220[255:0];
  _RAND_221 = {8{`RANDOM}};
  mem_221 = _RAND_221[255:0];
  _RAND_222 = {8{`RANDOM}};
  mem_222 = _RAND_222[255:0];
  _RAND_223 = {8{`RANDOM}};
  mem_223 = _RAND_223[255:0];
  _RAND_224 = {8{`RANDOM}};
  mem_224 = _RAND_224[255:0];
  _RAND_225 = {8{`RANDOM}};
  mem_225 = _RAND_225[255:0];
  _RAND_226 = {8{`RANDOM}};
  mem_226 = _RAND_226[255:0];
  _RAND_227 = {8{`RANDOM}};
  mem_227 = _RAND_227[255:0];
  _RAND_228 = {8{`RANDOM}};
  mem_228 = _RAND_228[255:0];
  _RAND_229 = {8{`RANDOM}};
  mem_229 = _RAND_229[255:0];
  _RAND_230 = {8{`RANDOM}};
  mem_230 = _RAND_230[255:0];
  _RAND_231 = {8{`RANDOM}};
  mem_231 = _RAND_231[255:0];
  _RAND_232 = {8{`RANDOM}};
  mem_232 = _RAND_232[255:0];
  _RAND_233 = {8{`RANDOM}};
  mem_233 = _RAND_233[255:0];
  _RAND_234 = {8{`RANDOM}};
  mem_234 = _RAND_234[255:0];
  _RAND_235 = {8{`RANDOM}};
  mem_235 = _RAND_235[255:0];
  _RAND_236 = {8{`RANDOM}};
  mem_236 = _RAND_236[255:0];
  _RAND_237 = {8{`RANDOM}};
  mem_237 = _RAND_237[255:0];
  _RAND_238 = {8{`RANDOM}};
  mem_238 = _RAND_238[255:0];
  _RAND_239 = {8{`RANDOM}};
  mem_239 = _RAND_239[255:0];
  _RAND_240 = {8{`RANDOM}};
  mem_240 = _RAND_240[255:0];
  _RAND_241 = {8{`RANDOM}};
  mem_241 = _RAND_241[255:0];
  _RAND_242 = {8{`RANDOM}};
  mem_242 = _RAND_242[255:0];
  _RAND_243 = {8{`RANDOM}};
  mem_243 = _RAND_243[255:0];
  _RAND_244 = {8{`RANDOM}};
  mem_244 = _RAND_244[255:0];
  _RAND_245 = {8{`RANDOM}};
  mem_245 = _RAND_245[255:0];
  _RAND_246 = {8{`RANDOM}};
  mem_246 = _RAND_246[255:0];
  _RAND_247 = {8{`RANDOM}};
  mem_247 = _RAND_247[255:0];
  _RAND_248 = {8{`RANDOM}};
  mem_248 = _RAND_248[255:0];
  _RAND_249 = {8{`RANDOM}};
  mem_249 = _RAND_249[255:0];
  _RAND_250 = {8{`RANDOM}};
  mem_250 = _RAND_250[255:0];
  _RAND_251 = {8{`RANDOM}};
  mem_251 = _RAND_251[255:0];
  _RAND_252 = {8{`RANDOM}};
  mem_252 = _RAND_252[255:0];
  _RAND_253 = {8{`RANDOM}};
  mem_253 = _RAND_253[255:0];
  _RAND_254 = {8{`RANDOM}};
  mem_254 = _RAND_254[255:0];
  _RAND_255 = {8{`RANDOM}};
  mem_255 = _RAND_255[255:0];
  _RAND_256 = {8{`RANDOM}};
  mem_256 = _RAND_256[255:0];
  _RAND_257 = {8{`RANDOM}};
  mem_257 = _RAND_257[255:0];
  _RAND_258 = {8{`RANDOM}};
  mem_258 = _RAND_258[255:0];
  _RAND_259 = {8{`RANDOM}};
  mem_259 = _RAND_259[255:0];
  _RAND_260 = {8{`RANDOM}};
  mem_260 = _RAND_260[255:0];
  _RAND_261 = {8{`RANDOM}};
  mem_261 = _RAND_261[255:0];
  _RAND_262 = {8{`RANDOM}};
  mem_262 = _RAND_262[255:0];
  _RAND_263 = {8{`RANDOM}};
  mem_263 = _RAND_263[255:0];
  _RAND_264 = {8{`RANDOM}};
  mem_264 = _RAND_264[255:0];
  _RAND_265 = {8{`RANDOM}};
  mem_265 = _RAND_265[255:0];
  _RAND_266 = {8{`RANDOM}};
  mem_266 = _RAND_266[255:0];
  _RAND_267 = {8{`RANDOM}};
  mem_267 = _RAND_267[255:0];
  _RAND_268 = {8{`RANDOM}};
  mem_268 = _RAND_268[255:0];
  _RAND_269 = {8{`RANDOM}};
  mem_269 = _RAND_269[255:0];
  _RAND_270 = {8{`RANDOM}};
  mem_270 = _RAND_270[255:0];
  _RAND_271 = {8{`RANDOM}};
  mem_271 = _RAND_271[255:0];
  _RAND_272 = {8{`RANDOM}};
  mem_272 = _RAND_272[255:0];
  _RAND_273 = {8{`RANDOM}};
  mem_273 = _RAND_273[255:0];
  _RAND_274 = {8{`RANDOM}};
  mem_274 = _RAND_274[255:0];
  _RAND_275 = {8{`RANDOM}};
  mem_275 = _RAND_275[255:0];
  _RAND_276 = {8{`RANDOM}};
  mem_276 = _RAND_276[255:0];
  _RAND_277 = {8{`RANDOM}};
  mem_277 = _RAND_277[255:0];
  _RAND_278 = {8{`RANDOM}};
  mem_278 = _RAND_278[255:0];
  _RAND_279 = {8{`RANDOM}};
  mem_279 = _RAND_279[255:0];
  _RAND_280 = {8{`RANDOM}};
  mem_280 = _RAND_280[255:0];
  _RAND_281 = {8{`RANDOM}};
  mem_281 = _RAND_281[255:0];
  _RAND_282 = {8{`RANDOM}};
  mem_282 = _RAND_282[255:0];
  _RAND_283 = {8{`RANDOM}};
  mem_283 = _RAND_283[255:0];
  _RAND_284 = {8{`RANDOM}};
  mem_284 = _RAND_284[255:0];
  _RAND_285 = {8{`RANDOM}};
  mem_285 = _RAND_285[255:0];
  _RAND_286 = {8{`RANDOM}};
  mem_286 = _RAND_286[255:0];
  _RAND_287 = {8{`RANDOM}};
  mem_287 = _RAND_287[255:0];
  _RAND_288 = {8{`RANDOM}};
  mem_288 = _RAND_288[255:0];
  _RAND_289 = {8{`RANDOM}};
  mem_289 = _RAND_289[255:0];
  _RAND_290 = {8{`RANDOM}};
  mem_290 = _RAND_290[255:0];
  _RAND_291 = {8{`RANDOM}};
  mem_291 = _RAND_291[255:0];
  _RAND_292 = {8{`RANDOM}};
  mem_292 = _RAND_292[255:0];
  _RAND_293 = {8{`RANDOM}};
  mem_293 = _RAND_293[255:0];
  _RAND_294 = {8{`RANDOM}};
  mem_294 = _RAND_294[255:0];
  _RAND_295 = {8{`RANDOM}};
  mem_295 = _RAND_295[255:0];
  _RAND_296 = {8{`RANDOM}};
  mem_296 = _RAND_296[255:0];
  _RAND_297 = {8{`RANDOM}};
  mem_297 = _RAND_297[255:0];
  _RAND_298 = {8{`RANDOM}};
  mem_298 = _RAND_298[255:0];
  _RAND_299 = {8{`RANDOM}};
  mem_299 = _RAND_299[255:0];
  _RAND_300 = {8{`RANDOM}};
  mem_300 = _RAND_300[255:0];
  _RAND_301 = {8{`RANDOM}};
  mem_301 = _RAND_301[255:0];
  _RAND_302 = {8{`RANDOM}};
  mem_302 = _RAND_302[255:0];
  _RAND_303 = {8{`RANDOM}};
  mem_303 = _RAND_303[255:0];
  _RAND_304 = {8{`RANDOM}};
  mem_304 = _RAND_304[255:0];
  _RAND_305 = {8{`RANDOM}};
  mem_305 = _RAND_305[255:0];
  _RAND_306 = {8{`RANDOM}};
  mem_306 = _RAND_306[255:0];
  _RAND_307 = {8{`RANDOM}};
  mem_307 = _RAND_307[255:0];
  _RAND_308 = {8{`RANDOM}};
  mem_308 = _RAND_308[255:0];
  _RAND_309 = {8{`RANDOM}};
  mem_309 = _RAND_309[255:0];
  _RAND_310 = {8{`RANDOM}};
  mem_310 = _RAND_310[255:0];
  _RAND_311 = {8{`RANDOM}};
  mem_311 = _RAND_311[255:0];
  _RAND_312 = {8{`RANDOM}};
  mem_312 = _RAND_312[255:0];
  _RAND_313 = {8{`RANDOM}};
  mem_313 = _RAND_313[255:0];
  _RAND_314 = {8{`RANDOM}};
  mem_314 = _RAND_314[255:0];
  _RAND_315 = {8{`RANDOM}};
  mem_315 = _RAND_315[255:0];
  _RAND_316 = {8{`RANDOM}};
  mem_316 = _RAND_316[255:0];
  _RAND_317 = {8{`RANDOM}};
  mem_317 = _RAND_317[255:0];
  _RAND_318 = {8{`RANDOM}};
  mem_318 = _RAND_318[255:0];
  _RAND_319 = {8{`RANDOM}};
  mem_319 = _RAND_319[255:0];
  _RAND_320 = {8{`RANDOM}};
  mem_320 = _RAND_320[255:0];
  _RAND_321 = {8{`RANDOM}};
  mem_321 = _RAND_321[255:0];
  _RAND_322 = {8{`RANDOM}};
  mem_322 = _RAND_322[255:0];
  _RAND_323 = {8{`RANDOM}};
  mem_323 = _RAND_323[255:0];
  _RAND_324 = {8{`RANDOM}};
  mem_324 = _RAND_324[255:0];
  _RAND_325 = {8{`RANDOM}};
  mem_325 = _RAND_325[255:0];
  _RAND_326 = {8{`RANDOM}};
  mem_326 = _RAND_326[255:0];
  _RAND_327 = {8{`RANDOM}};
  mem_327 = _RAND_327[255:0];
  _RAND_328 = {8{`RANDOM}};
  mem_328 = _RAND_328[255:0];
  _RAND_329 = {8{`RANDOM}};
  mem_329 = _RAND_329[255:0];
  _RAND_330 = {8{`RANDOM}};
  mem_330 = _RAND_330[255:0];
  _RAND_331 = {8{`RANDOM}};
  mem_331 = _RAND_331[255:0];
  _RAND_332 = {8{`RANDOM}};
  mem_332 = _RAND_332[255:0];
  _RAND_333 = {8{`RANDOM}};
  mem_333 = _RAND_333[255:0];
  _RAND_334 = {8{`RANDOM}};
  mem_334 = _RAND_334[255:0];
  _RAND_335 = {8{`RANDOM}};
  mem_335 = _RAND_335[255:0];
  _RAND_336 = {8{`RANDOM}};
  mem_336 = _RAND_336[255:0];
  _RAND_337 = {8{`RANDOM}};
  mem_337 = _RAND_337[255:0];
  _RAND_338 = {8{`RANDOM}};
  mem_338 = _RAND_338[255:0];
  _RAND_339 = {8{`RANDOM}};
  mem_339 = _RAND_339[255:0];
  _RAND_340 = {8{`RANDOM}};
  mem_340 = _RAND_340[255:0];
  _RAND_341 = {8{`RANDOM}};
  mem_341 = _RAND_341[255:0];
  _RAND_342 = {8{`RANDOM}};
  mem_342 = _RAND_342[255:0];
  _RAND_343 = {8{`RANDOM}};
  mem_343 = _RAND_343[255:0];
  _RAND_344 = {8{`RANDOM}};
  mem_344 = _RAND_344[255:0];
  _RAND_345 = {8{`RANDOM}};
  mem_345 = _RAND_345[255:0];
  _RAND_346 = {8{`RANDOM}};
  mem_346 = _RAND_346[255:0];
  _RAND_347 = {8{`RANDOM}};
  mem_347 = _RAND_347[255:0];
  _RAND_348 = {8{`RANDOM}};
  mem_348 = _RAND_348[255:0];
  _RAND_349 = {8{`RANDOM}};
  mem_349 = _RAND_349[255:0];
  _RAND_350 = {8{`RANDOM}};
  mem_350 = _RAND_350[255:0];
  _RAND_351 = {8{`RANDOM}};
  mem_351 = _RAND_351[255:0];
  _RAND_352 = {8{`RANDOM}};
  mem_352 = _RAND_352[255:0];
  _RAND_353 = {8{`RANDOM}};
  mem_353 = _RAND_353[255:0];
  _RAND_354 = {8{`RANDOM}};
  mem_354 = _RAND_354[255:0];
  _RAND_355 = {8{`RANDOM}};
  mem_355 = _RAND_355[255:0];
  _RAND_356 = {8{`RANDOM}};
  mem_356 = _RAND_356[255:0];
  _RAND_357 = {8{`RANDOM}};
  mem_357 = _RAND_357[255:0];
  _RAND_358 = {8{`RANDOM}};
  mem_358 = _RAND_358[255:0];
  _RAND_359 = {8{`RANDOM}};
  mem_359 = _RAND_359[255:0];
  _RAND_360 = {8{`RANDOM}};
  mem_360 = _RAND_360[255:0];
  _RAND_361 = {8{`RANDOM}};
  mem_361 = _RAND_361[255:0];
  _RAND_362 = {8{`RANDOM}};
  mem_362 = _RAND_362[255:0];
  _RAND_363 = {8{`RANDOM}};
  mem_363 = _RAND_363[255:0];
  _RAND_364 = {8{`RANDOM}};
  mem_364 = _RAND_364[255:0];
  _RAND_365 = {8{`RANDOM}};
  mem_365 = _RAND_365[255:0];
  _RAND_366 = {8{`RANDOM}};
  mem_366 = _RAND_366[255:0];
  _RAND_367 = {8{`RANDOM}};
  mem_367 = _RAND_367[255:0];
  _RAND_368 = {8{`RANDOM}};
  mem_368 = _RAND_368[255:0];
  _RAND_369 = {8{`RANDOM}};
  mem_369 = _RAND_369[255:0];
  _RAND_370 = {8{`RANDOM}};
  mem_370 = _RAND_370[255:0];
  _RAND_371 = {8{`RANDOM}};
  mem_371 = _RAND_371[255:0];
  _RAND_372 = {8{`RANDOM}};
  mem_372 = _RAND_372[255:0];
  _RAND_373 = {8{`RANDOM}};
  mem_373 = _RAND_373[255:0];
  _RAND_374 = {8{`RANDOM}};
  mem_374 = _RAND_374[255:0];
  _RAND_375 = {8{`RANDOM}};
  mem_375 = _RAND_375[255:0];
  _RAND_376 = {8{`RANDOM}};
  mem_376 = _RAND_376[255:0];
  _RAND_377 = {8{`RANDOM}};
  mem_377 = _RAND_377[255:0];
  _RAND_378 = {8{`RANDOM}};
  mem_378 = _RAND_378[255:0];
  _RAND_379 = {8{`RANDOM}};
  mem_379 = _RAND_379[255:0];
  _RAND_380 = {8{`RANDOM}};
  mem_380 = _RAND_380[255:0];
  _RAND_381 = {8{`RANDOM}};
  mem_381 = _RAND_381[255:0];
  _RAND_382 = {8{`RANDOM}};
  mem_382 = _RAND_382[255:0];
  _RAND_383 = {8{`RANDOM}};
  mem_383 = _RAND_383[255:0];
  _RAND_384 = {8{`RANDOM}};
  mem_384 = _RAND_384[255:0];
  _RAND_385 = {8{`RANDOM}};
  mem_385 = _RAND_385[255:0];
  _RAND_386 = {8{`RANDOM}};
  mem_386 = _RAND_386[255:0];
  _RAND_387 = {8{`RANDOM}};
  mem_387 = _RAND_387[255:0];
  _RAND_388 = {8{`RANDOM}};
  mem_388 = _RAND_388[255:0];
  _RAND_389 = {8{`RANDOM}};
  mem_389 = _RAND_389[255:0];
  _RAND_390 = {8{`RANDOM}};
  mem_390 = _RAND_390[255:0];
  _RAND_391 = {8{`RANDOM}};
  mem_391 = _RAND_391[255:0];
  _RAND_392 = {8{`RANDOM}};
  mem_392 = _RAND_392[255:0];
  _RAND_393 = {8{`RANDOM}};
  mem_393 = _RAND_393[255:0];
  _RAND_394 = {8{`RANDOM}};
  mem_394 = _RAND_394[255:0];
  _RAND_395 = {8{`RANDOM}};
  mem_395 = _RAND_395[255:0];
  _RAND_396 = {8{`RANDOM}};
  mem_396 = _RAND_396[255:0];
  _RAND_397 = {8{`RANDOM}};
  mem_397 = _RAND_397[255:0];
  _RAND_398 = {8{`RANDOM}};
  mem_398 = _RAND_398[255:0];
  _RAND_399 = {8{`RANDOM}};
  mem_399 = _RAND_399[255:0];
  _RAND_400 = {8{`RANDOM}};
  mem_400 = _RAND_400[255:0];
  _RAND_401 = {8{`RANDOM}};
  mem_401 = _RAND_401[255:0];
  _RAND_402 = {8{`RANDOM}};
  mem_402 = _RAND_402[255:0];
  _RAND_403 = {8{`RANDOM}};
  mem_403 = _RAND_403[255:0];
  _RAND_404 = {8{`RANDOM}};
  mem_404 = _RAND_404[255:0];
  _RAND_405 = {8{`RANDOM}};
  mem_405 = _RAND_405[255:0];
  _RAND_406 = {8{`RANDOM}};
  mem_406 = _RAND_406[255:0];
  _RAND_407 = {8{`RANDOM}};
  mem_407 = _RAND_407[255:0];
  _RAND_408 = {8{`RANDOM}};
  mem_408 = _RAND_408[255:0];
  _RAND_409 = {8{`RANDOM}};
  mem_409 = _RAND_409[255:0];
  _RAND_410 = {8{`RANDOM}};
  mem_410 = _RAND_410[255:0];
  _RAND_411 = {8{`RANDOM}};
  mem_411 = _RAND_411[255:0];
  _RAND_412 = {8{`RANDOM}};
  mem_412 = _RAND_412[255:0];
  _RAND_413 = {8{`RANDOM}};
  mem_413 = _RAND_413[255:0];
  _RAND_414 = {8{`RANDOM}};
  mem_414 = _RAND_414[255:0];
  _RAND_415 = {8{`RANDOM}};
  mem_415 = _RAND_415[255:0];
  _RAND_416 = {8{`RANDOM}};
  mem_416 = _RAND_416[255:0];
  _RAND_417 = {8{`RANDOM}};
  mem_417 = _RAND_417[255:0];
  _RAND_418 = {8{`RANDOM}};
  mem_418 = _RAND_418[255:0];
  _RAND_419 = {8{`RANDOM}};
  mem_419 = _RAND_419[255:0];
  _RAND_420 = {8{`RANDOM}};
  mem_420 = _RAND_420[255:0];
  _RAND_421 = {8{`RANDOM}};
  mem_421 = _RAND_421[255:0];
  _RAND_422 = {8{`RANDOM}};
  mem_422 = _RAND_422[255:0];
  _RAND_423 = {8{`RANDOM}};
  mem_423 = _RAND_423[255:0];
  _RAND_424 = {8{`RANDOM}};
  mem_424 = _RAND_424[255:0];
  _RAND_425 = {8{`RANDOM}};
  mem_425 = _RAND_425[255:0];
  _RAND_426 = {8{`RANDOM}};
  mem_426 = _RAND_426[255:0];
  _RAND_427 = {8{`RANDOM}};
  mem_427 = _RAND_427[255:0];
  _RAND_428 = {8{`RANDOM}};
  mem_428 = _RAND_428[255:0];
  _RAND_429 = {8{`RANDOM}};
  mem_429 = _RAND_429[255:0];
  _RAND_430 = {8{`RANDOM}};
  mem_430 = _RAND_430[255:0];
  _RAND_431 = {8{`RANDOM}};
  mem_431 = _RAND_431[255:0];
  _RAND_432 = {8{`RANDOM}};
  mem_432 = _RAND_432[255:0];
  _RAND_433 = {8{`RANDOM}};
  mem_433 = _RAND_433[255:0];
  _RAND_434 = {8{`RANDOM}};
  mem_434 = _RAND_434[255:0];
  _RAND_435 = {8{`RANDOM}};
  mem_435 = _RAND_435[255:0];
  _RAND_436 = {8{`RANDOM}};
  mem_436 = _RAND_436[255:0];
  _RAND_437 = {8{`RANDOM}};
  mem_437 = _RAND_437[255:0];
  _RAND_438 = {8{`RANDOM}};
  mem_438 = _RAND_438[255:0];
  _RAND_439 = {8{`RANDOM}};
  mem_439 = _RAND_439[255:0];
  _RAND_440 = {8{`RANDOM}};
  mem_440 = _RAND_440[255:0];
  _RAND_441 = {8{`RANDOM}};
  mem_441 = _RAND_441[255:0];
  _RAND_442 = {8{`RANDOM}};
  mem_442 = _RAND_442[255:0];
  _RAND_443 = {8{`RANDOM}};
  mem_443 = _RAND_443[255:0];
  _RAND_444 = {8{`RANDOM}};
  mem_444 = _RAND_444[255:0];
  _RAND_445 = {8{`RANDOM}};
  mem_445 = _RAND_445[255:0];
  _RAND_446 = {8{`RANDOM}};
  mem_446 = _RAND_446[255:0];
  _RAND_447 = {8{`RANDOM}};
  mem_447 = _RAND_447[255:0];
  _RAND_448 = {8{`RANDOM}};
  mem_448 = _RAND_448[255:0];
  _RAND_449 = {8{`RANDOM}};
  mem_449 = _RAND_449[255:0];
  _RAND_450 = {8{`RANDOM}};
  mem_450 = _RAND_450[255:0];
  _RAND_451 = {8{`RANDOM}};
  mem_451 = _RAND_451[255:0];
  _RAND_452 = {8{`RANDOM}};
  mem_452 = _RAND_452[255:0];
  _RAND_453 = {8{`RANDOM}};
  mem_453 = _RAND_453[255:0];
  _RAND_454 = {8{`RANDOM}};
  mem_454 = _RAND_454[255:0];
  _RAND_455 = {8{`RANDOM}};
  mem_455 = _RAND_455[255:0];
  _RAND_456 = {8{`RANDOM}};
  mem_456 = _RAND_456[255:0];
  _RAND_457 = {8{`RANDOM}};
  mem_457 = _RAND_457[255:0];
  _RAND_458 = {8{`RANDOM}};
  mem_458 = _RAND_458[255:0];
  _RAND_459 = {8{`RANDOM}};
  mem_459 = _RAND_459[255:0];
  _RAND_460 = {8{`RANDOM}};
  mem_460 = _RAND_460[255:0];
  _RAND_461 = {8{`RANDOM}};
  mem_461 = _RAND_461[255:0];
  _RAND_462 = {8{`RANDOM}};
  mem_462 = _RAND_462[255:0];
  _RAND_463 = {8{`RANDOM}};
  mem_463 = _RAND_463[255:0];
  _RAND_464 = {8{`RANDOM}};
  mem_464 = _RAND_464[255:0];
  _RAND_465 = {8{`RANDOM}};
  mem_465 = _RAND_465[255:0];
  _RAND_466 = {8{`RANDOM}};
  mem_466 = _RAND_466[255:0];
  _RAND_467 = {8{`RANDOM}};
  mem_467 = _RAND_467[255:0];
  _RAND_468 = {8{`RANDOM}};
  mem_468 = _RAND_468[255:0];
  _RAND_469 = {8{`RANDOM}};
  mem_469 = _RAND_469[255:0];
  _RAND_470 = {8{`RANDOM}};
  mem_470 = _RAND_470[255:0];
  _RAND_471 = {8{`RANDOM}};
  mem_471 = _RAND_471[255:0];
  _RAND_472 = {8{`RANDOM}};
  mem_472 = _RAND_472[255:0];
  _RAND_473 = {8{`RANDOM}};
  mem_473 = _RAND_473[255:0];
  _RAND_474 = {8{`RANDOM}};
  mem_474 = _RAND_474[255:0];
  _RAND_475 = {8{`RANDOM}};
  mem_475 = _RAND_475[255:0];
  _RAND_476 = {8{`RANDOM}};
  mem_476 = _RAND_476[255:0];
  _RAND_477 = {8{`RANDOM}};
  mem_477 = _RAND_477[255:0];
  _RAND_478 = {8{`RANDOM}};
  mem_478 = _RAND_478[255:0];
  _RAND_479 = {8{`RANDOM}};
  mem_479 = _RAND_479[255:0];
  _RAND_480 = {8{`RANDOM}};
  mem_480 = _RAND_480[255:0];
  _RAND_481 = {8{`RANDOM}};
  mem_481 = _RAND_481[255:0];
  _RAND_482 = {8{`RANDOM}};
  mem_482 = _RAND_482[255:0];
  _RAND_483 = {8{`RANDOM}};
  mem_483 = _RAND_483[255:0];
  _RAND_484 = {8{`RANDOM}};
  mem_484 = _RAND_484[255:0];
  _RAND_485 = {8{`RANDOM}};
  mem_485 = _RAND_485[255:0];
  _RAND_486 = {8{`RANDOM}};
  mem_486 = _RAND_486[255:0];
  _RAND_487 = {8{`RANDOM}};
  mem_487 = _RAND_487[255:0];
  _RAND_488 = {8{`RANDOM}};
  mem_488 = _RAND_488[255:0];
  _RAND_489 = {8{`RANDOM}};
  mem_489 = _RAND_489[255:0];
  _RAND_490 = {8{`RANDOM}};
  mem_490 = _RAND_490[255:0];
  _RAND_491 = {8{`RANDOM}};
  mem_491 = _RAND_491[255:0];
  _RAND_492 = {8{`RANDOM}};
  mem_492 = _RAND_492[255:0];
  _RAND_493 = {8{`RANDOM}};
  mem_493 = _RAND_493[255:0];
  _RAND_494 = {8{`RANDOM}};
  mem_494 = _RAND_494[255:0];
  _RAND_495 = {8{`RANDOM}};
  mem_495 = _RAND_495[255:0];
  _RAND_496 = {8{`RANDOM}};
  mem_496 = _RAND_496[255:0];
  _RAND_497 = {8{`RANDOM}};
  mem_497 = _RAND_497[255:0];
  _RAND_498 = {8{`RANDOM}};
  mem_498 = _RAND_498[255:0];
  _RAND_499 = {8{`RANDOM}};
  mem_499 = _RAND_499[255:0];
  _RAND_500 = {8{`RANDOM}};
  mem_500 = _RAND_500[255:0];
  _RAND_501 = {8{`RANDOM}};
  mem_501 = _RAND_501[255:0];
  _RAND_502 = {8{`RANDOM}};
  mem_502 = _RAND_502[255:0];
  _RAND_503 = {8{`RANDOM}};
  mem_503 = _RAND_503[255:0];
  _RAND_504 = {8{`RANDOM}};
  mem_504 = _RAND_504[255:0];
  _RAND_505 = {8{`RANDOM}};
  mem_505 = _RAND_505[255:0];
  _RAND_506 = {8{`RANDOM}};
  mem_506 = _RAND_506[255:0];
  _RAND_507 = {8{`RANDOM}};
  mem_507 = _RAND_507[255:0];
  _RAND_508 = {8{`RANDOM}};
  mem_508 = _RAND_508[255:0];
  _RAND_509 = {8{`RANDOM}};
  mem_509 = _RAND_509[255:0];
  _RAND_510 = {8{`RANDOM}};
  mem_510 = _RAND_510[255:0];
  _RAND_511 = {8{`RANDOM}};
  mem_511 = _RAND_511[255:0];
  _RAND_512 = {8{`RANDOM}};
  io_douta_REG = _RAND_512[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM_2(
  input          clock,
  input          reset,
  input          io_web,
  input  [8:0]   io_addra,
  input  [8:0]   io_addrb,
  input  [255:0] io_dinb,
  output [255:0] io_douta
);
  wire  sim_dual_port_bram_clock; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_reset; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_io_web; // @[RAMWrapper.scala 30:36]
  wire [8:0] sim_dual_port_bram_io_addra; // @[RAMWrapper.scala 30:36]
  wire [8:0] sim_dual_port_bram_io_addrb; // @[RAMWrapper.scala 30:36]
  wire [255:0] sim_dual_port_bram_io_dinb; // @[RAMWrapper.scala 30:36]
  wire [255:0] sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 30:36]
  SimDualPortBRAM_2 sim_dual_port_bram ( // @[RAMWrapper.scala 30:36]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_web(sim_dual_port_bram_io_web),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dinb(sim_dual_port_bram_io_dinb),
    .io_douta(sim_dual_port_bram_io_douta)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_web = io_web; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_dinb = io_dinb; // @[RAMWrapper.scala 31:27]
endmodule
module SimDualPortBRAM_3(
  input         clock,
  input         reset,
  input         io_web,
  input  [8:0]  io_addra,
  input  [8:0]  io_addrb,
  input  [19:0] io_dinb,
  output [19:0] io_douta
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem_0; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_1; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_2; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_3; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_4; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_5; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_6; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_7; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_8; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_9; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_10; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_11; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_12; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_13; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_14; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_15; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_16; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_17; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_18; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_19; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_20; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_21; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_22; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_23; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_24; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_25; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_26; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_27; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_28; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_29; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_30; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_31; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_32; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_33; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_34; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_35; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_36; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_37; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_38; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_39; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_40; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_41; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_42; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_43; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_44; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_45; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_46; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_47; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_48; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_49; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_50; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_51; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_52; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_53; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_54; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_55; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_56; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_57; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_58; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_59; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_60; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_61; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_62; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_63; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_64; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_65; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_66; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_67; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_68; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_69; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_70; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_71; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_72; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_73; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_74; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_75; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_76; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_77; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_78; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_79; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_80; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_81; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_82; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_83; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_84; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_85; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_86; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_87; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_88; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_89; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_90; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_91; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_92; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_93; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_94; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_95; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_96; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_97; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_98; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_99; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_100; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_101; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_102; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_103; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_104; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_105; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_106; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_107; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_108; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_109; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_110; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_111; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_112; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_113; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_114; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_115; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_116; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_117; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_118; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_119; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_120; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_121; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_122; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_123; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_124; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_125; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_126; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_127; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_128; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_129; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_130; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_131; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_132; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_133; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_134; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_135; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_136; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_137; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_138; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_139; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_140; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_141; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_142; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_143; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_144; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_145; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_146; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_147; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_148; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_149; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_150; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_151; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_152; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_153; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_154; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_155; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_156; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_157; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_158; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_159; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_160; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_161; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_162; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_163; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_164; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_165; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_166; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_167; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_168; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_169; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_170; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_171; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_172; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_173; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_174; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_175; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_176; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_177; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_178; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_179; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_180; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_181; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_182; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_183; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_184; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_185; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_186; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_187; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_188; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_189; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_190; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_191; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_192; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_193; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_194; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_195; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_196; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_197; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_198; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_199; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_200; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_201; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_202; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_203; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_204; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_205; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_206; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_207; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_208; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_209; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_210; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_211; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_212; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_213; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_214; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_215; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_216; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_217; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_218; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_219; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_220; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_221; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_222; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_223; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_224; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_225; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_226; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_227; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_228; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_229; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_230; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_231; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_232; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_233; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_234; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_235; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_236; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_237; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_238; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_239; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_240; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_241; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_242; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_243; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_244; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_245; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_246; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_247; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_248; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_249; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_250; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_251; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_252; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_253; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_254; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_255; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_256; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_257; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_258; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_259; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_260; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_261; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_262; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_263; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_264; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_265; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_266; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_267; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_268; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_269; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_270; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_271; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_272; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_273; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_274; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_275; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_276; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_277; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_278; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_279; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_280; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_281; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_282; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_283; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_284; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_285; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_286; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_287; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_288; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_289; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_290; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_291; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_292; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_293; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_294; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_295; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_296; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_297; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_298; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_299; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_300; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_301; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_302; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_303; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_304; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_305; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_306; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_307; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_308; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_309; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_310; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_311; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_312; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_313; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_314; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_315; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_316; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_317; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_318; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_319; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_320; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_321; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_322; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_323; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_324; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_325; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_326; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_327; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_328; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_329; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_330; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_331; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_332; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_333; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_334; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_335; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_336; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_337; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_338; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_339; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_340; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_341; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_342; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_343; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_344; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_345; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_346; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_347; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_348; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_349; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_350; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_351; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_352; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_353; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_354; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_355; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_356; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_357; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_358; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_359; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_360; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_361; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_362; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_363; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_364; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_365; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_366; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_367; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_368; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_369; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_370; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_371; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_372; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_373; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_374; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_375; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_376; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_377; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_378; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_379; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_380; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_381; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_382; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_383; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_384; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_385; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_386; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_387; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_388; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_389; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_390; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_391; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_392; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_393; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_394; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_395; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_396; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_397; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_398; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_399; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_400; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_401; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_402; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_403; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_404; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_405; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_406; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_407; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_408; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_409; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_410; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_411; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_412; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_413; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_414; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_415; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_416; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_417; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_418; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_419; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_420; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_421; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_422; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_423; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_424; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_425; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_426; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_427; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_428; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_429; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_430; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_431; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_432; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_433; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_434; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_435; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_436; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_437; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_438; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_439; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_440; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_441; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_442; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_443; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_444; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_445; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_446; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_447; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_448; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_449; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_450; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_451; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_452; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_453; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_454; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_455; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_456; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_457; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_458; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_459; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_460; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_461; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_462; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_463; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_464; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_465; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_466; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_467; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_468; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_469; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_470; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_471; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_472; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_473; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_474; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_475; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_476; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_477; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_478; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_479; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_480; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_481; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_482; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_483; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_484; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_485; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_486; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_487; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_488; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_489; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_490; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_491; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_492; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_493; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_494; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_495; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_496; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_497; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_498; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_499; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_500; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_501; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_502; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_503; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_504; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_505; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_506; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_507; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_508; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_509; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_510; // @[RAMWrapper.scala 41:20]
  reg [19:0] mem_511; // @[RAMWrapper.scala 41:20]
  reg [19:0] io_douta_REG; // @[RAMWrapper.scala 43:22]
  wire [19:0] _GEN_1 = 9'h1 == io_addra ? mem_1 : mem_0; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_2 = 9'h2 == io_addra ? mem_2 : _GEN_1; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_3 = 9'h3 == io_addra ? mem_3 : _GEN_2; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_4 = 9'h4 == io_addra ? mem_4 : _GEN_3; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_5 = 9'h5 == io_addra ? mem_5 : _GEN_4; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_6 = 9'h6 == io_addra ? mem_6 : _GEN_5; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_7 = 9'h7 == io_addra ? mem_7 : _GEN_6; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_8 = 9'h8 == io_addra ? mem_8 : _GEN_7; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_9 = 9'h9 == io_addra ? mem_9 : _GEN_8; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_10 = 9'ha == io_addra ? mem_10 : _GEN_9; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_11 = 9'hb == io_addra ? mem_11 : _GEN_10; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_12 = 9'hc == io_addra ? mem_12 : _GEN_11; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_13 = 9'hd == io_addra ? mem_13 : _GEN_12; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_14 = 9'he == io_addra ? mem_14 : _GEN_13; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_15 = 9'hf == io_addra ? mem_15 : _GEN_14; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_16 = 9'h10 == io_addra ? mem_16 : _GEN_15; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_17 = 9'h11 == io_addra ? mem_17 : _GEN_16; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_18 = 9'h12 == io_addra ? mem_18 : _GEN_17; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_19 = 9'h13 == io_addra ? mem_19 : _GEN_18; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_20 = 9'h14 == io_addra ? mem_20 : _GEN_19; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_21 = 9'h15 == io_addra ? mem_21 : _GEN_20; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_22 = 9'h16 == io_addra ? mem_22 : _GEN_21; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_23 = 9'h17 == io_addra ? mem_23 : _GEN_22; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_24 = 9'h18 == io_addra ? mem_24 : _GEN_23; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_25 = 9'h19 == io_addra ? mem_25 : _GEN_24; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_26 = 9'h1a == io_addra ? mem_26 : _GEN_25; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_27 = 9'h1b == io_addra ? mem_27 : _GEN_26; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_28 = 9'h1c == io_addra ? mem_28 : _GEN_27; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_29 = 9'h1d == io_addra ? mem_29 : _GEN_28; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_30 = 9'h1e == io_addra ? mem_30 : _GEN_29; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_31 = 9'h1f == io_addra ? mem_31 : _GEN_30; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_32 = 9'h20 == io_addra ? mem_32 : _GEN_31; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_33 = 9'h21 == io_addra ? mem_33 : _GEN_32; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_34 = 9'h22 == io_addra ? mem_34 : _GEN_33; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_35 = 9'h23 == io_addra ? mem_35 : _GEN_34; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_36 = 9'h24 == io_addra ? mem_36 : _GEN_35; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_37 = 9'h25 == io_addra ? mem_37 : _GEN_36; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_38 = 9'h26 == io_addra ? mem_38 : _GEN_37; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_39 = 9'h27 == io_addra ? mem_39 : _GEN_38; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_40 = 9'h28 == io_addra ? mem_40 : _GEN_39; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_41 = 9'h29 == io_addra ? mem_41 : _GEN_40; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_42 = 9'h2a == io_addra ? mem_42 : _GEN_41; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_43 = 9'h2b == io_addra ? mem_43 : _GEN_42; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_44 = 9'h2c == io_addra ? mem_44 : _GEN_43; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_45 = 9'h2d == io_addra ? mem_45 : _GEN_44; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_46 = 9'h2e == io_addra ? mem_46 : _GEN_45; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_47 = 9'h2f == io_addra ? mem_47 : _GEN_46; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_48 = 9'h30 == io_addra ? mem_48 : _GEN_47; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_49 = 9'h31 == io_addra ? mem_49 : _GEN_48; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_50 = 9'h32 == io_addra ? mem_50 : _GEN_49; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_51 = 9'h33 == io_addra ? mem_51 : _GEN_50; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_52 = 9'h34 == io_addra ? mem_52 : _GEN_51; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_53 = 9'h35 == io_addra ? mem_53 : _GEN_52; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_54 = 9'h36 == io_addra ? mem_54 : _GEN_53; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_55 = 9'h37 == io_addra ? mem_55 : _GEN_54; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_56 = 9'h38 == io_addra ? mem_56 : _GEN_55; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_57 = 9'h39 == io_addra ? mem_57 : _GEN_56; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_58 = 9'h3a == io_addra ? mem_58 : _GEN_57; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_59 = 9'h3b == io_addra ? mem_59 : _GEN_58; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_60 = 9'h3c == io_addra ? mem_60 : _GEN_59; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_61 = 9'h3d == io_addra ? mem_61 : _GEN_60; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_62 = 9'h3e == io_addra ? mem_62 : _GEN_61; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_63 = 9'h3f == io_addra ? mem_63 : _GEN_62; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_64 = 9'h40 == io_addra ? mem_64 : _GEN_63; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_65 = 9'h41 == io_addra ? mem_65 : _GEN_64; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_66 = 9'h42 == io_addra ? mem_66 : _GEN_65; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_67 = 9'h43 == io_addra ? mem_67 : _GEN_66; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_68 = 9'h44 == io_addra ? mem_68 : _GEN_67; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_69 = 9'h45 == io_addra ? mem_69 : _GEN_68; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_70 = 9'h46 == io_addra ? mem_70 : _GEN_69; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_71 = 9'h47 == io_addra ? mem_71 : _GEN_70; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_72 = 9'h48 == io_addra ? mem_72 : _GEN_71; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_73 = 9'h49 == io_addra ? mem_73 : _GEN_72; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_74 = 9'h4a == io_addra ? mem_74 : _GEN_73; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_75 = 9'h4b == io_addra ? mem_75 : _GEN_74; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_76 = 9'h4c == io_addra ? mem_76 : _GEN_75; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_77 = 9'h4d == io_addra ? mem_77 : _GEN_76; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_78 = 9'h4e == io_addra ? mem_78 : _GEN_77; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_79 = 9'h4f == io_addra ? mem_79 : _GEN_78; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_80 = 9'h50 == io_addra ? mem_80 : _GEN_79; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_81 = 9'h51 == io_addra ? mem_81 : _GEN_80; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_82 = 9'h52 == io_addra ? mem_82 : _GEN_81; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_83 = 9'h53 == io_addra ? mem_83 : _GEN_82; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_84 = 9'h54 == io_addra ? mem_84 : _GEN_83; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_85 = 9'h55 == io_addra ? mem_85 : _GEN_84; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_86 = 9'h56 == io_addra ? mem_86 : _GEN_85; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_87 = 9'h57 == io_addra ? mem_87 : _GEN_86; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_88 = 9'h58 == io_addra ? mem_88 : _GEN_87; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_89 = 9'h59 == io_addra ? mem_89 : _GEN_88; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_90 = 9'h5a == io_addra ? mem_90 : _GEN_89; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_91 = 9'h5b == io_addra ? mem_91 : _GEN_90; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_92 = 9'h5c == io_addra ? mem_92 : _GEN_91; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_93 = 9'h5d == io_addra ? mem_93 : _GEN_92; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_94 = 9'h5e == io_addra ? mem_94 : _GEN_93; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_95 = 9'h5f == io_addra ? mem_95 : _GEN_94; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_96 = 9'h60 == io_addra ? mem_96 : _GEN_95; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_97 = 9'h61 == io_addra ? mem_97 : _GEN_96; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_98 = 9'h62 == io_addra ? mem_98 : _GEN_97; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_99 = 9'h63 == io_addra ? mem_99 : _GEN_98; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_100 = 9'h64 == io_addra ? mem_100 : _GEN_99; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_101 = 9'h65 == io_addra ? mem_101 : _GEN_100; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_102 = 9'h66 == io_addra ? mem_102 : _GEN_101; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_103 = 9'h67 == io_addra ? mem_103 : _GEN_102; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_104 = 9'h68 == io_addra ? mem_104 : _GEN_103; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_105 = 9'h69 == io_addra ? mem_105 : _GEN_104; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_106 = 9'h6a == io_addra ? mem_106 : _GEN_105; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_107 = 9'h6b == io_addra ? mem_107 : _GEN_106; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_108 = 9'h6c == io_addra ? mem_108 : _GEN_107; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_109 = 9'h6d == io_addra ? mem_109 : _GEN_108; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_110 = 9'h6e == io_addra ? mem_110 : _GEN_109; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_111 = 9'h6f == io_addra ? mem_111 : _GEN_110; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_112 = 9'h70 == io_addra ? mem_112 : _GEN_111; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_113 = 9'h71 == io_addra ? mem_113 : _GEN_112; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_114 = 9'h72 == io_addra ? mem_114 : _GEN_113; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_115 = 9'h73 == io_addra ? mem_115 : _GEN_114; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_116 = 9'h74 == io_addra ? mem_116 : _GEN_115; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_117 = 9'h75 == io_addra ? mem_117 : _GEN_116; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_118 = 9'h76 == io_addra ? mem_118 : _GEN_117; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_119 = 9'h77 == io_addra ? mem_119 : _GEN_118; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_120 = 9'h78 == io_addra ? mem_120 : _GEN_119; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_121 = 9'h79 == io_addra ? mem_121 : _GEN_120; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_122 = 9'h7a == io_addra ? mem_122 : _GEN_121; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_123 = 9'h7b == io_addra ? mem_123 : _GEN_122; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_124 = 9'h7c == io_addra ? mem_124 : _GEN_123; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_125 = 9'h7d == io_addra ? mem_125 : _GEN_124; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_126 = 9'h7e == io_addra ? mem_126 : _GEN_125; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_127 = 9'h7f == io_addra ? mem_127 : _GEN_126; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_128 = 9'h80 == io_addra ? mem_128 : _GEN_127; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_129 = 9'h81 == io_addra ? mem_129 : _GEN_128; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_130 = 9'h82 == io_addra ? mem_130 : _GEN_129; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_131 = 9'h83 == io_addra ? mem_131 : _GEN_130; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_132 = 9'h84 == io_addra ? mem_132 : _GEN_131; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_133 = 9'h85 == io_addra ? mem_133 : _GEN_132; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_134 = 9'h86 == io_addra ? mem_134 : _GEN_133; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_135 = 9'h87 == io_addra ? mem_135 : _GEN_134; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_136 = 9'h88 == io_addra ? mem_136 : _GEN_135; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_137 = 9'h89 == io_addra ? mem_137 : _GEN_136; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_138 = 9'h8a == io_addra ? mem_138 : _GEN_137; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_139 = 9'h8b == io_addra ? mem_139 : _GEN_138; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_140 = 9'h8c == io_addra ? mem_140 : _GEN_139; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_141 = 9'h8d == io_addra ? mem_141 : _GEN_140; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_142 = 9'h8e == io_addra ? mem_142 : _GEN_141; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_143 = 9'h8f == io_addra ? mem_143 : _GEN_142; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_144 = 9'h90 == io_addra ? mem_144 : _GEN_143; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_145 = 9'h91 == io_addra ? mem_145 : _GEN_144; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_146 = 9'h92 == io_addra ? mem_146 : _GEN_145; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_147 = 9'h93 == io_addra ? mem_147 : _GEN_146; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_148 = 9'h94 == io_addra ? mem_148 : _GEN_147; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_149 = 9'h95 == io_addra ? mem_149 : _GEN_148; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_150 = 9'h96 == io_addra ? mem_150 : _GEN_149; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_151 = 9'h97 == io_addra ? mem_151 : _GEN_150; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_152 = 9'h98 == io_addra ? mem_152 : _GEN_151; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_153 = 9'h99 == io_addra ? mem_153 : _GEN_152; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_154 = 9'h9a == io_addra ? mem_154 : _GEN_153; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_155 = 9'h9b == io_addra ? mem_155 : _GEN_154; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_156 = 9'h9c == io_addra ? mem_156 : _GEN_155; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_157 = 9'h9d == io_addra ? mem_157 : _GEN_156; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_158 = 9'h9e == io_addra ? mem_158 : _GEN_157; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_159 = 9'h9f == io_addra ? mem_159 : _GEN_158; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_160 = 9'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_161 = 9'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_162 = 9'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_163 = 9'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_164 = 9'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_165 = 9'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_166 = 9'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_167 = 9'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_168 = 9'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_169 = 9'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_170 = 9'haa == io_addra ? mem_170 : _GEN_169; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_171 = 9'hab == io_addra ? mem_171 : _GEN_170; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_172 = 9'hac == io_addra ? mem_172 : _GEN_171; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_173 = 9'had == io_addra ? mem_173 : _GEN_172; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_174 = 9'hae == io_addra ? mem_174 : _GEN_173; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_175 = 9'haf == io_addra ? mem_175 : _GEN_174; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_176 = 9'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_177 = 9'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_178 = 9'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_179 = 9'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_180 = 9'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_181 = 9'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_182 = 9'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_183 = 9'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_184 = 9'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_185 = 9'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_186 = 9'hba == io_addra ? mem_186 : _GEN_185; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_187 = 9'hbb == io_addra ? mem_187 : _GEN_186; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_188 = 9'hbc == io_addra ? mem_188 : _GEN_187; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_189 = 9'hbd == io_addra ? mem_189 : _GEN_188; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_190 = 9'hbe == io_addra ? mem_190 : _GEN_189; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_191 = 9'hbf == io_addra ? mem_191 : _GEN_190; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_192 = 9'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_193 = 9'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_194 = 9'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_195 = 9'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_196 = 9'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_197 = 9'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_198 = 9'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_199 = 9'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_200 = 9'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_201 = 9'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_202 = 9'hca == io_addra ? mem_202 : _GEN_201; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_203 = 9'hcb == io_addra ? mem_203 : _GEN_202; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_204 = 9'hcc == io_addra ? mem_204 : _GEN_203; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_205 = 9'hcd == io_addra ? mem_205 : _GEN_204; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_206 = 9'hce == io_addra ? mem_206 : _GEN_205; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_207 = 9'hcf == io_addra ? mem_207 : _GEN_206; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_208 = 9'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_209 = 9'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_210 = 9'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_211 = 9'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_212 = 9'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_213 = 9'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_214 = 9'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_215 = 9'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_216 = 9'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_217 = 9'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_218 = 9'hda == io_addra ? mem_218 : _GEN_217; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_219 = 9'hdb == io_addra ? mem_219 : _GEN_218; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_220 = 9'hdc == io_addra ? mem_220 : _GEN_219; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_221 = 9'hdd == io_addra ? mem_221 : _GEN_220; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_222 = 9'hde == io_addra ? mem_222 : _GEN_221; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_223 = 9'hdf == io_addra ? mem_223 : _GEN_222; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_224 = 9'he0 == io_addra ? mem_224 : _GEN_223; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_225 = 9'he1 == io_addra ? mem_225 : _GEN_224; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_226 = 9'he2 == io_addra ? mem_226 : _GEN_225; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_227 = 9'he3 == io_addra ? mem_227 : _GEN_226; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_228 = 9'he4 == io_addra ? mem_228 : _GEN_227; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_229 = 9'he5 == io_addra ? mem_229 : _GEN_228; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_230 = 9'he6 == io_addra ? mem_230 : _GEN_229; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_231 = 9'he7 == io_addra ? mem_231 : _GEN_230; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_232 = 9'he8 == io_addra ? mem_232 : _GEN_231; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_233 = 9'he9 == io_addra ? mem_233 : _GEN_232; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_234 = 9'hea == io_addra ? mem_234 : _GEN_233; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_235 = 9'heb == io_addra ? mem_235 : _GEN_234; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_236 = 9'hec == io_addra ? mem_236 : _GEN_235; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_237 = 9'hed == io_addra ? mem_237 : _GEN_236; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_238 = 9'hee == io_addra ? mem_238 : _GEN_237; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_239 = 9'hef == io_addra ? mem_239 : _GEN_238; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_240 = 9'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_241 = 9'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_242 = 9'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_243 = 9'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_244 = 9'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_245 = 9'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_246 = 9'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_247 = 9'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_248 = 9'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_249 = 9'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_250 = 9'hfa == io_addra ? mem_250 : _GEN_249; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_251 = 9'hfb == io_addra ? mem_251 : _GEN_250; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_252 = 9'hfc == io_addra ? mem_252 : _GEN_251; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_253 = 9'hfd == io_addra ? mem_253 : _GEN_252; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_254 = 9'hfe == io_addra ? mem_254 : _GEN_253; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_255 = 9'hff == io_addra ? mem_255 : _GEN_254; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_256 = 9'h100 == io_addra ? mem_256 : _GEN_255; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_257 = 9'h101 == io_addra ? mem_257 : _GEN_256; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_258 = 9'h102 == io_addra ? mem_258 : _GEN_257; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_259 = 9'h103 == io_addra ? mem_259 : _GEN_258; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_260 = 9'h104 == io_addra ? mem_260 : _GEN_259; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_261 = 9'h105 == io_addra ? mem_261 : _GEN_260; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_262 = 9'h106 == io_addra ? mem_262 : _GEN_261; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_263 = 9'h107 == io_addra ? mem_263 : _GEN_262; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_264 = 9'h108 == io_addra ? mem_264 : _GEN_263; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_265 = 9'h109 == io_addra ? mem_265 : _GEN_264; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_266 = 9'h10a == io_addra ? mem_266 : _GEN_265; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_267 = 9'h10b == io_addra ? mem_267 : _GEN_266; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_268 = 9'h10c == io_addra ? mem_268 : _GEN_267; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_269 = 9'h10d == io_addra ? mem_269 : _GEN_268; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_270 = 9'h10e == io_addra ? mem_270 : _GEN_269; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_271 = 9'h10f == io_addra ? mem_271 : _GEN_270; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_272 = 9'h110 == io_addra ? mem_272 : _GEN_271; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_273 = 9'h111 == io_addra ? mem_273 : _GEN_272; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_274 = 9'h112 == io_addra ? mem_274 : _GEN_273; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_275 = 9'h113 == io_addra ? mem_275 : _GEN_274; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_276 = 9'h114 == io_addra ? mem_276 : _GEN_275; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_277 = 9'h115 == io_addra ? mem_277 : _GEN_276; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_278 = 9'h116 == io_addra ? mem_278 : _GEN_277; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_279 = 9'h117 == io_addra ? mem_279 : _GEN_278; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_280 = 9'h118 == io_addra ? mem_280 : _GEN_279; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_281 = 9'h119 == io_addra ? mem_281 : _GEN_280; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_282 = 9'h11a == io_addra ? mem_282 : _GEN_281; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_283 = 9'h11b == io_addra ? mem_283 : _GEN_282; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_284 = 9'h11c == io_addra ? mem_284 : _GEN_283; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_285 = 9'h11d == io_addra ? mem_285 : _GEN_284; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_286 = 9'h11e == io_addra ? mem_286 : _GEN_285; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_287 = 9'h11f == io_addra ? mem_287 : _GEN_286; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_288 = 9'h120 == io_addra ? mem_288 : _GEN_287; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_289 = 9'h121 == io_addra ? mem_289 : _GEN_288; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_290 = 9'h122 == io_addra ? mem_290 : _GEN_289; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_291 = 9'h123 == io_addra ? mem_291 : _GEN_290; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_292 = 9'h124 == io_addra ? mem_292 : _GEN_291; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_293 = 9'h125 == io_addra ? mem_293 : _GEN_292; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_294 = 9'h126 == io_addra ? mem_294 : _GEN_293; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_295 = 9'h127 == io_addra ? mem_295 : _GEN_294; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_296 = 9'h128 == io_addra ? mem_296 : _GEN_295; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_297 = 9'h129 == io_addra ? mem_297 : _GEN_296; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_298 = 9'h12a == io_addra ? mem_298 : _GEN_297; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_299 = 9'h12b == io_addra ? mem_299 : _GEN_298; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_300 = 9'h12c == io_addra ? mem_300 : _GEN_299; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_301 = 9'h12d == io_addra ? mem_301 : _GEN_300; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_302 = 9'h12e == io_addra ? mem_302 : _GEN_301; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_303 = 9'h12f == io_addra ? mem_303 : _GEN_302; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_304 = 9'h130 == io_addra ? mem_304 : _GEN_303; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_305 = 9'h131 == io_addra ? mem_305 : _GEN_304; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_306 = 9'h132 == io_addra ? mem_306 : _GEN_305; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_307 = 9'h133 == io_addra ? mem_307 : _GEN_306; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_308 = 9'h134 == io_addra ? mem_308 : _GEN_307; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_309 = 9'h135 == io_addra ? mem_309 : _GEN_308; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_310 = 9'h136 == io_addra ? mem_310 : _GEN_309; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_311 = 9'h137 == io_addra ? mem_311 : _GEN_310; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_312 = 9'h138 == io_addra ? mem_312 : _GEN_311; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_313 = 9'h139 == io_addra ? mem_313 : _GEN_312; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_314 = 9'h13a == io_addra ? mem_314 : _GEN_313; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_315 = 9'h13b == io_addra ? mem_315 : _GEN_314; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_316 = 9'h13c == io_addra ? mem_316 : _GEN_315; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_317 = 9'h13d == io_addra ? mem_317 : _GEN_316; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_318 = 9'h13e == io_addra ? mem_318 : _GEN_317; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_319 = 9'h13f == io_addra ? mem_319 : _GEN_318; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_320 = 9'h140 == io_addra ? mem_320 : _GEN_319; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_321 = 9'h141 == io_addra ? mem_321 : _GEN_320; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_322 = 9'h142 == io_addra ? mem_322 : _GEN_321; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_323 = 9'h143 == io_addra ? mem_323 : _GEN_322; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_324 = 9'h144 == io_addra ? mem_324 : _GEN_323; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_325 = 9'h145 == io_addra ? mem_325 : _GEN_324; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_326 = 9'h146 == io_addra ? mem_326 : _GEN_325; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_327 = 9'h147 == io_addra ? mem_327 : _GEN_326; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_328 = 9'h148 == io_addra ? mem_328 : _GEN_327; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_329 = 9'h149 == io_addra ? mem_329 : _GEN_328; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_330 = 9'h14a == io_addra ? mem_330 : _GEN_329; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_331 = 9'h14b == io_addra ? mem_331 : _GEN_330; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_332 = 9'h14c == io_addra ? mem_332 : _GEN_331; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_333 = 9'h14d == io_addra ? mem_333 : _GEN_332; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_334 = 9'h14e == io_addra ? mem_334 : _GEN_333; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_335 = 9'h14f == io_addra ? mem_335 : _GEN_334; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_336 = 9'h150 == io_addra ? mem_336 : _GEN_335; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_337 = 9'h151 == io_addra ? mem_337 : _GEN_336; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_338 = 9'h152 == io_addra ? mem_338 : _GEN_337; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_339 = 9'h153 == io_addra ? mem_339 : _GEN_338; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_340 = 9'h154 == io_addra ? mem_340 : _GEN_339; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_341 = 9'h155 == io_addra ? mem_341 : _GEN_340; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_342 = 9'h156 == io_addra ? mem_342 : _GEN_341; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_343 = 9'h157 == io_addra ? mem_343 : _GEN_342; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_344 = 9'h158 == io_addra ? mem_344 : _GEN_343; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_345 = 9'h159 == io_addra ? mem_345 : _GEN_344; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_346 = 9'h15a == io_addra ? mem_346 : _GEN_345; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_347 = 9'h15b == io_addra ? mem_347 : _GEN_346; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_348 = 9'h15c == io_addra ? mem_348 : _GEN_347; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_349 = 9'h15d == io_addra ? mem_349 : _GEN_348; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_350 = 9'h15e == io_addra ? mem_350 : _GEN_349; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_351 = 9'h15f == io_addra ? mem_351 : _GEN_350; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_352 = 9'h160 == io_addra ? mem_352 : _GEN_351; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_353 = 9'h161 == io_addra ? mem_353 : _GEN_352; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_354 = 9'h162 == io_addra ? mem_354 : _GEN_353; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_355 = 9'h163 == io_addra ? mem_355 : _GEN_354; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_356 = 9'h164 == io_addra ? mem_356 : _GEN_355; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_357 = 9'h165 == io_addra ? mem_357 : _GEN_356; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_358 = 9'h166 == io_addra ? mem_358 : _GEN_357; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_359 = 9'h167 == io_addra ? mem_359 : _GEN_358; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_360 = 9'h168 == io_addra ? mem_360 : _GEN_359; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_361 = 9'h169 == io_addra ? mem_361 : _GEN_360; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_362 = 9'h16a == io_addra ? mem_362 : _GEN_361; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_363 = 9'h16b == io_addra ? mem_363 : _GEN_362; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_364 = 9'h16c == io_addra ? mem_364 : _GEN_363; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_365 = 9'h16d == io_addra ? mem_365 : _GEN_364; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_366 = 9'h16e == io_addra ? mem_366 : _GEN_365; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_367 = 9'h16f == io_addra ? mem_367 : _GEN_366; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_368 = 9'h170 == io_addra ? mem_368 : _GEN_367; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_369 = 9'h171 == io_addra ? mem_369 : _GEN_368; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_370 = 9'h172 == io_addra ? mem_370 : _GEN_369; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_371 = 9'h173 == io_addra ? mem_371 : _GEN_370; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_372 = 9'h174 == io_addra ? mem_372 : _GEN_371; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_373 = 9'h175 == io_addra ? mem_373 : _GEN_372; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_374 = 9'h176 == io_addra ? mem_374 : _GEN_373; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_375 = 9'h177 == io_addra ? mem_375 : _GEN_374; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_376 = 9'h178 == io_addra ? mem_376 : _GEN_375; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_377 = 9'h179 == io_addra ? mem_377 : _GEN_376; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_378 = 9'h17a == io_addra ? mem_378 : _GEN_377; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_379 = 9'h17b == io_addra ? mem_379 : _GEN_378; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_380 = 9'h17c == io_addra ? mem_380 : _GEN_379; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_381 = 9'h17d == io_addra ? mem_381 : _GEN_380; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_382 = 9'h17e == io_addra ? mem_382 : _GEN_381; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_383 = 9'h17f == io_addra ? mem_383 : _GEN_382; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_384 = 9'h180 == io_addra ? mem_384 : _GEN_383; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_385 = 9'h181 == io_addra ? mem_385 : _GEN_384; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_386 = 9'h182 == io_addra ? mem_386 : _GEN_385; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_387 = 9'h183 == io_addra ? mem_387 : _GEN_386; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_388 = 9'h184 == io_addra ? mem_388 : _GEN_387; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_389 = 9'h185 == io_addra ? mem_389 : _GEN_388; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_390 = 9'h186 == io_addra ? mem_390 : _GEN_389; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_391 = 9'h187 == io_addra ? mem_391 : _GEN_390; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_392 = 9'h188 == io_addra ? mem_392 : _GEN_391; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_393 = 9'h189 == io_addra ? mem_393 : _GEN_392; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_394 = 9'h18a == io_addra ? mem_394 : _GEN_393; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_395 = 9'h18b == io_addra ? mem_395 : _GEN_394; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_396 = 9'h18c == io_addra ? mem_396 : _GEN_395; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_397 = 9'h18d == io_addra ? mem_397 : _GEN_396; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_398 = 9'h18e == io_addra ? mem_398 : _GEN_397; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_399 = 9'h18f == io_addra ? mem_399 : _GEN_398; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_400 = 9'h190 == io_addra ? mem_400 : _GEN_399; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_401 = 9'h191 == io_addra ? mem_401 : _GEN_400; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_402 = 9'h192 == io_addra ? mem_402 : _GEN_401; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_403 = 9'h193 == io_addra ? mem_403 : _GEN_402; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_404 = 9'h194 == io_addra ? mem_404 : _GEN_403; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_405 = 9'h195 == io_addra ? mem_405 : _GEN_404; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_406 = 9'h196 == io_addra ? mem_406 : _GEN_405; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_407 = 9'h197 == io_addra ? mem_407 : _GEN_406; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_408 = 9'h198 == io_addra ? mem_408 : _GEN_407; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_409 = 9'h199 == io_addra ? mem_409 : _GEN_408; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_410 = 9'h19a == io_addra ? mem_410 : _GEN_409; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_411 = 9'h19b == io_addra ? mem_411 : _GEN_410; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_412 = 9'h19c == io_addra ? mem_412 : _GEN_411; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_413 = 9'h19d == io_addra ? mem_413 : _GEN_412; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_414 = 9'h19e == io_addra ? mem_414 : _GEN_413; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_415 = 9'h19f == io_addra ? mem_415 : _GEN_414; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_416 = 9'h1a0 == io_addra ? mem_416 : _GEN_415; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_417 = 9'h1a1 == io_addra ? mem_417 : _GEN_416; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_418 = 9'h1a2 == io_addra ? mem_418 : _GEN_417; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_419 = 9'h1a3 == io_addra ? mem_419 : _GEN_418; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_420 = 9'h1a4 == io_addra ? mem_420 : _GEN_419; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_421 = 9'h1a5 == io_addra ? mem_421 : _GEN_420; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_422 = 9'h1a6 == io_addra ? mem_422 : _GEN_421; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_423 = 9'h1a7 == io_addra ? mem_423 : _GEN_422; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_424 = 9'h1a8 == io_addra ? mem_424 : _GEN_423; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_425 = 9'h1a9 == io_addra ? mem_425 : _GEN_424; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_426 = 9'h1aa == io_addra ? mem_426 : _GEN_425; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_427 = 9'h1ab == io_addra ? mem_427 : _GEN_426; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_428 = 9'h1ac == io_addra ? mem_428 : _GEN_427; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_429 = 9'h1ad == io_addra ? mem_429 : _GEN_428; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_430 = 9'h1ae == io_addra ? mem_430 : _GEN_429; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_431 = 9'h1af == io_addra ? mem_431 : _GEN_430; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_432 = 9'h1b0 == io_addra ? mem_432 : _GEN_431; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_433 = 9'h1b1 == io_addra ? mem_433 : _GEN_432; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_434 = 9'h1b2 == io_addra ? mem_434 : _GEN_433; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_435 = 9'h1b3 == io_addra ? mem_435 : _GEN_434; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_436 = 9'h1b4 == io_addra ? mem_436 : _GEN_435; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_437 = 9'h1b5 == io_addra ? mem_437 : _GEN_436; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_438 = 9'h1b6 == io_addra ? mem_438 : _GEN_437; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_439 = 9'h1b7 == io_addra ? mem_439 : _GEN_438; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_440 = 9'h1b8 == io_addra ? mem_440 : _GEN_439; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_441 = 9'h1b9 == io_addra ? mem_441 : _GEN_440; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_442 = 9'h1ba == io_addra ? mem_442 : _GEN_441; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_443 = 9'h1bb == io_addra ? mem_443 : _GEN_442; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_444 = 9'h1bc == io_addra ? mem_444 : _GEN_443; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_445 = 9'h1bd == io_addra ? mem_445 : _GEN_444; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_446 = 9'h1be == io_addra ? mem_446 : _GEN_445; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_447 = 9'h1bf == io_addra ? mem_447 : _GEN_446; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_448 = 9'h1c0 == io_addra ? mem_448 : _GEN_447; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_449 = 9'h1c1 == io_addra ? mem_449 : _GEN_448; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_450 = 9'h1c2 == io_addra ? mem_450 : _GEN_449; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_451 = 9'h1c3 == io_addra ? mem_451 : _GEN_450; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_452 = 9'h1c4 == io_addra ? mem_452 : _GEN_451; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_453 = 9'h1c5 == io_addra ? mem_453 : _GEN_452; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_454 = 9'h1c6 == io_addra ? mem_454 : _GEN_453; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_455 = 9'h1c7 == io_addra ? mem_455 : _GEN_454; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_456 = 9'h1c8 == io_addra ? mem_456 : _GEN_455; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_457 = 9'h1c9 == io_addra ? mem_457 : _GEN_456; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_458 = 9'h1ca == io_addra ? mem_458 : _GEN_457; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_459 = 9'h1cb == io_addra ? mem_459 : _GEN_458; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_460 = 9'h1cc == io_addra ? mem_460 : _GEN_459; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_461 = 9'h1cd == io_addra ? mem_461 : _GEN_460; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_462 = 9'h1ce == io_addra ? mem_462 : _GEN_461; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_463 = 9'h1cf == io_addra ? mem_463 : _GEN_462; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_464 = 9'h1d0 == io_addra ? mem_464 : _GEN_463; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_465 = 9'h1d1 == io_addra ? mem_465 : _GEN_464; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_466 = 9'h1d2 == io_addra ? mem_466 : _GEN_465; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_467 = 9'h1d3 == io_addra ? mem_467 : _GEN_466; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_468 = 9'h1d4 == io_addra ? mem_468 : _GEN_467; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_469 = 9'h1d5 == io_addra ? mem_469 : _GEN_468; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_470 = 9'h1d6 == io_addra ? mem_470 : _GEN_469; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_471 = 9'h1d7 == io_addra ? mem_471 : _GEN_470; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_472 = 9'h1d8 == io_addra ? mem_472 : _GEN_471; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_473 = 9'h1d9 == io_addra ? mem_473 : _GEN_472; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_474 = 9'h1da == io_addra ? mem_474 : _GEN_473; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_475 = 9'h1db == io_addra ? mem_475 : _GEN_474; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_476 = 9'h1dc == io_addra ? mem_476 : _GEN_475; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_477 = 9'h1dd == io_addra ? mem_477 : _GEN_476; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_478 = 9'h1de == io_addra ? mem_478 : _GEN_477; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_479 = 9'h1df == io_addra ? mem_479 : _GEN_478; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_480 = 9'h1e0 == io_addra ? mem_480 : _GEN_479; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_481 = 9'h1e1 == io_addra ? mem_481 : _GEN_480; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_482 = 9'h1e2 == io_addra ? mem_482 : _GEN_481; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_483 = 9'h1e3 == io_addra ? mem_483 : _GEN_482; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_484 = 9'h1e4 == io_addra ? mem_484 : _GEN_483; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_485 = 9'h1e5 == io_addra ? mem_485 : _GEN_484; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_486 = 9'h1e6 == io_addra ? mem_486 : _GEN_485; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_487 = 9'h1e7 == io_addra ? mem_487 : _GEN_486; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_488 = 9'h1e8 == io_addra ? mem_488 : _GEN_487; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_489 = 9'h1e9 == io_addra ? mem_489 : _GEN_488; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_490 = 9'h1ea == io_addra ? mem_490 : _GEN_489; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_491 = 9'h1eb == io_addra ? mem_491 : _GEN_490; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_492 = 9'h1ec == io_addra ? mem_492 : _GEN_491; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_493 = 9'h1ed == io_addra ? mem_493 : _GEN_492; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_494 = 9'h1ee == io_addra ? mem_494 : _GEN_493; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_495 = 9'h1ef == io_addra ? mem_495 : _GEN_494; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_496 = 9'h1f0 == io_addra ? mem_496 : _GEN_495; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_497 = 9'h1f1 == io_addra ? mem_497 : _GEN_496; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_498 = 9'h1f2 == io_addra ? mem_498 : _GEN_497; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_499 = 9'h1f3 == io_addra ? mem_499 : _GEN_498; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_500 = 9'h1f4 == io_addra ? mem_500 : _GEN_499; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_501 = 9'h1f5 == io_addra ? mem_501 : _GEN_500; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_502 = 9'h1f6 == io_addra ? mem_502 : _GEN_501; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_503 = 9'h1f7 == io_addra ? mem_503 : _GEN_502; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_504 = 9'h1f8 == io_addra ? mem_504 : _GEN_503; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_505 = 9'h1f9 == io_addra ? mem_505 : _GEN_504; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_506 = 9'h1fa == io_addra ? mem_506 : _GEN_505; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  wire [19:0] _GEN_507 = 9'h1fb == io_addra ? mem_507 : _GEN_506; // @[RAMWrapper.scala 43:22 RAMWrapper.scala 43:22]
  assign io_douta = io_douta_REG; // @[RAMWrapper.scala 43:12]
  always @(posedge clock) begin
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_0 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_0 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_1 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_1 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_2 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_2 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_3 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_3 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_4 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_4 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_5 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_5 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_6 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_6 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_7 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_7 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_8 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_8 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_9 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_9 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_10 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_10 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_11 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_11 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_12 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_12 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_13 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_13 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_14 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_14 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_15 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_15 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_16 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_16 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_17 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_17 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_18 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_18 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_19 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_19 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_20 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_20 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_21 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_21 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_22 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_22 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_23 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_23 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_24 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_24 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_25 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_25 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_26 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_26 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_27 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_27 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_28 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_28 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_29 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_29 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_30 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_30 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_31 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_31 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_32 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h20 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_32 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_33 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h21 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_33 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_34 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h22 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_34 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_35 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h23 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_35 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_36 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h24 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_36 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_37 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h25 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_37 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_38 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h26 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_38 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_39 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h27 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_39 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_40 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h28 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_40 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_41 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h29 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_41 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_42 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_42 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_43 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_43 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_44 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_44 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_45 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_45 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_46 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_46 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_47 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h2f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_47 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_48 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h30 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_48 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_49 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h31 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_49 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_50 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h32 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_50 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_51 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h33 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_51 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_52 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h34 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_52 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_53 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h35 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_53 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_54 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h36 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_54 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_55 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h37 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_55 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_56 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h38 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_56 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_57 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h39 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_57 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_58 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_58 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_59 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_59 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_60 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_60 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_61 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_61 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_62 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_62 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_63 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h3f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_63 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_64 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h40 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_64 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_65 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h41 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_65 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_66 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h42 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_66 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_67 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h43 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_67 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_68 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h44 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_68 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_69 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h45 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_69 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_70 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h46 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_70 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_71 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h47 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_71 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_72 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h48 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_72 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_73 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h49 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_73 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_74 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_74 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_75 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_75 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_76 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_76 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_77 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_77 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_78 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_78 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_79 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h4f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_79 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_80 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h50 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_80 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_81 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h51 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_81 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_82 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h52 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_82 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_83 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h53 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_83 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_84 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h54 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_84 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_85 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h55 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_85 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_86 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h56 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_86 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_87 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h57 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_87 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_88 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h58 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_88 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_89 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h59 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_89 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_90 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_90 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_91 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_91 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_92 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_92 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_93 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_93 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_94 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_94 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_95 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h5f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_95 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_96 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h60 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_96 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_97 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h61 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_97 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_98 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h62 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_98 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_99 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h63 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_99 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_100 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h64 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_100 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_101 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h65 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_101 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_102 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h66 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_102 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_103 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h67 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_103 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_104 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h68 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_104 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_105 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h69 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_105 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_106 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_106 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_107 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_107 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_108 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_108 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_109 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_109 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_110 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_110 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_111 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h6f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_111 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_112 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h70 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_112 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_113 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h71 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_113 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_114 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h72 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_114 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_115 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h73 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_115 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_116 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h74 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_116 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_117 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h75 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_117 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_118 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h76 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_118 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_119 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h77 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_119 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_120 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h78 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_120 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_121 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h79 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_121 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_122 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_122 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_123 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_123 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_124 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_124 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_125 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_125 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_126 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_126 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_127 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h7f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_127 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_128 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h80 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_128 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_129 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h81 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_129 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_130 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h82 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_130 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_131 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h83 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_131 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_132 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h84 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_132 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_133 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h85 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_133 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_134 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h86 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_134 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_135 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h87 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_135 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_136 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h88 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_136 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_137 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h89 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_137 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_138 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_138 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_139 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_139 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_140 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_140 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_141 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_141 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_142 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_142 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_143 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h8f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_143 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_144 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h90 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_144 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_145 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h91 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_145 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_146 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h92 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_146 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_147 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h93 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_147 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_148 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h94 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_148 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_149 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h95 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_149 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_150 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h96 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_150 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_151 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h97 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_151 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_152 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h98 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_152 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_153 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h99 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_153 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_154 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_154 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_155 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_155 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_156 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_156 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_157 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_157 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_158 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_158 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_159 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h9f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_159 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_160 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_160 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_161 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_161 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_162 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_162 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_163 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_163 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_164 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_164 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_165 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_165 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_166 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_166 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_167 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_167 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_168 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_168 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_169 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'ha9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_169 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_170 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'haa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_170 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_171 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hab == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_171 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_172 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hac == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_172 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_173 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'had == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_173 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_174 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hae == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_174 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_175 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'haf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_175 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_176 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_176 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_177 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_177 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_178 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_178 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_179 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_179 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_180 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_180 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_181 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_181 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_182 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_182 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_183 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_183 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_184 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_184 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_185 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hb9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_185 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_186 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hba == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_186 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_187 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_187 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_188 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_188 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_189 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_189 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_190 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_190 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_191 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hbf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_191 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_192 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_192 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_193 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_193 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_194 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_194 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_195 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_195 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_196 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_196 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_197 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_197 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_198 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_198 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_199 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_199 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_200 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_200 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_201 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hc9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_201 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_202 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hca == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_202 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_203 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_203 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_204 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_204 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_205 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_205 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_206 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hce == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_206 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_207 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hcf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_207 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_208 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_208 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_209 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_209 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_210 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_210 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_211 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_211 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_212 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_212 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_213 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_213 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_214 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_214 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_215 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_215 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_216 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_216 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_217 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hd9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_217 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_218 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hda == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_218 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_219 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_219 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_220 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_220 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_221 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_221 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_222 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hde == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_222 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_223 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hdf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_223 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_224 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_224 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_225 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_225 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_226 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_226 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_227 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_227 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_228 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_228 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_229 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_229 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_230 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_230 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_231 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_231 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_232 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_232 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_233 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'he9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_233 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_234 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hea == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_234 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_235 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'heb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_235 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_236 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hec == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_236 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_237 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hed == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_237 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_238 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hee == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_238 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_239 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hef == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_239 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_240 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_240 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_241 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_241 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_242 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_242 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_243 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_243 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_244 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_244 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_245 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_245 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_246 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_246 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_247 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_247 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_248 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_248 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_249 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hf9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_249 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_250 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_250 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_251 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_251 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_252 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_252 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_253 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_253 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_254 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hfe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_254 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_255 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'hff == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_255 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_256 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h100 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_256 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_257 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h101 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_257 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_258 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h102 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_258 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_259 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h103 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_259 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_260 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h104 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_260 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_261 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h105 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_261 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_262 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h106 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_262 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_263 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h107 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_263 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_264 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h108 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_264 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_265 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h109 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_265 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_266 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_266 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_267 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_267 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_268 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_268 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_269 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_269 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_270 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_270 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_271 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h10f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_271 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_272 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h110 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_272 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_273 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h111 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_273 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_274 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h112 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_274 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_275 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h113 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_275 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_276 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h114 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_276 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_277 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h115 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_277 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_278 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h116 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_278 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_279 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h117 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_279 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_280 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h118 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_280 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_281 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h119 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_281 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_282 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_282 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_283 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_283 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_284 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_284 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_285 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_285 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_286 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_286 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_287 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h11f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_287 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_288 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h120 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_288 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_289 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h121 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_289 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_290 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h122 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_290 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_291 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h123 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_291 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_292 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h124 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_292 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_293 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h125 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_293 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_294 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h126 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_294 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_295 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h127 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_295 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_296 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h128 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_296 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_297 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h129 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_297 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_298 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_298 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_299 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_299 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_300 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_300 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_301 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_301 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_302 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_302 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_303 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h12f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_303 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_304 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h130 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_304 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_305 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h131 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_305 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_306 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h132 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_306 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_307 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h133 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_307 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_308 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h134 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_308 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_309 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h135 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_309 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_310 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h136 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_310 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_311 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h137 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_311 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_312 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h138 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_312 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_313 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h139 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_313 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_314 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_314 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_315 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_315 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_316 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_316 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_317 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_317 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_318 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_318 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_319 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h13f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_319 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_320 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h140 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_320 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_321 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h141 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_321 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_322 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h142 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_322 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_323 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h143 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_323 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_324 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h144 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_324 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_325 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h145 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_325 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_326 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h146 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_326 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_327 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h147 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_327 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_328 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h148 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_328 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_329 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h149 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_329 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_330 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_330 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_331 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_331 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_332 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_332 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_333 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_333 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_334 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_334 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_335 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h14f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_335 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_336 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h150 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_336 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_337 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h151 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_337 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_338 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h152 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_338 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_339 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h153 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_339 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_340 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h154 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_340 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_341 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h155 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_341 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_342 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h156 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_342 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_343 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h157 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_343 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_344 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h158 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_344 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_345 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h159 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_345 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_346 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_346 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_347 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_347 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_348 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_348 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_349 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_349 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_350 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_350 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_351 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h15f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_351 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_352 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h160 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_352 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_353 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h161 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_353 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_354 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h162 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_354 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_355 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h163 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_355 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_356 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h164 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_356 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_357 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h165 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_357 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_358 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h166 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_358 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_359 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h167 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_359 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_360 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h168 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_360 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_361 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h169 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_361 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_362 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_362 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_363 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_363 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_364 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_364 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_365 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_365 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_366 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_366 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_367 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h16f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_367 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_368 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h170 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_368 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_369 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h171 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_369 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_370 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h172 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_370 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_371 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h173 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_371 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_372 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h174 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_372 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_373 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h175 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_373 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_374 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h176 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_374 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_375 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h177 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_375 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_376 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h178 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_376 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_377 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h179 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_377 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_378 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_378 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_379 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_379 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_380 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_380 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_381 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_381 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_382 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_382 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_383 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h17f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_383 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_384 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h180 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_384 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_385 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h181 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_385 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_386 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h182 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_386 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_387 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h183 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_387 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_388 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h184 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_388 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_389 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h185 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_389 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_390 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h186 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_390 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_391 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h187 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_391 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_392 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h188 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_392 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_393 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h189 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_393 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_394 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_394 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_395 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_395 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_396 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_396 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_397 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_397 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_398 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_398 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_399 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h18f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_399 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_400 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h190 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_400 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_401 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h191 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_401 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_402 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h192 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_402 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_403 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h193 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_403 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_404 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h194 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_404 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_405 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h195 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_405 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_406 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h196 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_406 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_407 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h197 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_407 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_408 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h198 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_408 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_409 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h199 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_409 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_410 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19a == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_410 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_411 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19b == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_411 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_412 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19c == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_412 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_413 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19d == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_413 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_414 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19e == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_414 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_415 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h19f == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_415 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_416 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_416 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_417 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_417 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_418 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_418 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_419 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_419 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_420 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_420 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_421 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_421 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_422 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_422 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_423 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_423 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_424 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_424 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_425 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1a9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_425 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_426 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1aa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_426 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_427 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ab == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_427 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_428 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ac == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_428 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_429 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ad == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_429 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_430 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ae == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_430 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_431 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1af == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_431 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_432 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_432 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_433 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_433 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_434 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_434 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_435 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_435 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_436 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_436 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_437 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_437 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_438 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_438 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_439 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_439 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_440 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_440 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_441 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1b9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_441 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_442 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ba == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_442 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_443 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_443 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_444 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_444 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_445 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_445 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_446 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1be == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_446 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_447 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1bf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_447 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_448 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_448 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_449 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_449 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_450 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_450 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_451 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_451 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_452 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_452 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_453 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_453 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_454 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_454 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_455 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_455 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_456 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_456 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_457 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1c9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_457 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_458 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ca == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_458 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_459 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_459 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_460 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_460 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_461 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_461 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_462 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ce == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_462 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_463 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1cf == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_463 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_464 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_464 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_465 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_465 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_466 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_466 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_467 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_467 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_468 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_468 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_469 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_469 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_470 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_470 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_471 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_471 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_472 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_472 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_473 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1d9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_473 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_474 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1da == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_474 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_475 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1db == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_475 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_476 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1dc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_476 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_477 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1dd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_477 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_478 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1de == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_478 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_479 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1df == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_479 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_480 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_480 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_481 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_481 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_482 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_482 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_483 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_483 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_484 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_484 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_485 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_485 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_486 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_486 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_487 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_487 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_488 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_488 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_489 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1e9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_489 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_490 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ea == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_490 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_491 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1eb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_491 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_492 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ec == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_492 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_493 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ed == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_493 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_494 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ee == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_494 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_495 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ef == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_495 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_496 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f0 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_496 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_497 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f1 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_497 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_498 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f2 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_498 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_499 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f3 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_499 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_500 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f4 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_500 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_501 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f5 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_501 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_502 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f6 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_502 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_503 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f7 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_503 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_504 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f8 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_504 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_505 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1f9 == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_505 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_506 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fa == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_506 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_507 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fb == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_507 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_508 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fc == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_508 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_509 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fd == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_509 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_510 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1fe == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_510 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (reset) begin // @[RAMWrapper.scala 41:20]
      mem_511 <= 20'h0; // @[RAMWrapper.scala 41:20]
    end else if (io_web) begin // @[RAMWrapper.scala 49:16]
      if (9'h1ff == io_addrb) begin // @[RAMWrapper.scala 50:19]
        mem_511 <= io_dinb; // @[RAMWrapper.scala 50:19]
      end
    end
    if (9'h1ff == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_511; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fe == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_510; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fd == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_509; // @[RAMWrapper.scala 43:22]
    end else if (9'h1fc == io_addra) begin // @[RAMWrapper.scala 43:22]
      io_douta_REG <= mem_508; // @[RAMWrapper.scala 43:22]
    end else begin
      io_douta_REG <= _GEN_507;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[19:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[19:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[19:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[19:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[19:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[19:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[19:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[19:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[19:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[19:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[19:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[19:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[19:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[19:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[19:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[19:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[19:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[19:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[19:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[19:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[19:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[19:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[19:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[19:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[19:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[19:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[19:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[19:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[19:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[19:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[19:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[19:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[19:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[19:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[19:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[19:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[19:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[19:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[19:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[19:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[19:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[19:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[19:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[19:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[19:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[19:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[19:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[19:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[19:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[19:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[19:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[19:0];
  _RAND_128 = {1{`RANDOM}};
  mem_128 = _RAND_128[19:0];
  _RAND_129 = {1{`RANDOM}};
  mem_129 = _RAND_129[19:0];
  _RAND_130 = {1{`RANDOM}};
  mem_130 = _RAND_130[19:0];
  _RAND_131 = {1{`RANDOM}};
  mem_131 = _RAND_131[19:0];
  _RAND_132 = {1{`RANDOM}};
  mem_132 = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  mem_133 = _RAND_133[19:0];
  _RAND_134 = {1{`RANDOM}};
  mem_134 = _RAND_134[19:0];
  _RAND_135 = {1{`RANDOM}};
  mem_135 = _RAND_135[19:0];
  _RAND_136 = {1{`RANDOM}};
  mem_136 = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  mem_137 = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  mem_138 = _RAND_138[19:0];
  _RAND_139 = {1{`RANDOM}};
  mem_139 = _RAND_139[19:0];
  _RAND_140 = {1{`RANDOM}};
  mem_140 = _RAND_140[19:0];
  _RAND_141 = {1{`RANDOM}};
  mem_141 = _RAND_141[19:0];
  _RAND_142 = {1{`RANDOM}};
  mem_142 = _RAND_142[19:0];
  _RAND_143 = {1{`RANDOM}};
  mem_143 = _RAND_143[19:0];
  _RAND_144 = {1{`RANDOM}};
  mem_144 = _RAND_144[19:0];
  _RAND_145 = {1{`RANDOM}};
  mem_145 = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  mem_146 = _RAND_146[19:0];
  _RAND_147 = {1{`RANDOM}};
  mem_147 = _RAND_147[19:0];
  _RAND_148 = {1{`RANDOM}};
  mem_148 = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  mem_149 = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  mem_150 = _RAND_150[19:0];
  _RAND_151 = {1{`RANDOM}};
  mem_151 = _RAND_151[19:0];
  _RAND_152 = {1{`RANDOM}};
  mem_152 = _RAND_152[19:0];
  _RAND_153 = {1{`RANDOM}};
  mem_153 = _RAND_153[19:0];
  _RAND_154 = {1{`RANDOM}};
  mem_154 = _RAND_154[19:0];
  _RAND_155 = {1{`RANDOM}};
  mem_155 = _RAND_155[19:0];
  _RAND_156 = {1{`RANDOM}};
  mem_156 = _RAND_156[19:0];
  _RAND_157 = {1{`RANDOM}};
  mem_157 = _RAND_157[19:0];
  _RAND_158 = {1{`RANDOM}};
  mem_158 = _RAND_158[19:0];
  _RAND_159 = {1{`RANDOM}};
  mem_159 = _RAND_159[19:0];
  _RAND_160 = {1{`RANDOM}};
  mem_160 = _RAND_160[19:0];
  _RAND_161 = {1{`RANDOM}};
  mem_161 = _RAND_161[19:0];
  _RAND_162 = {1{`RANDOM}};
  mem_162 = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  mem_163 = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  mem_164 = _RAND_164[19:0];
  _RAND_165 = {1{`RANDOM}};
  mem_165 = _RAND_165[19:0];
  _RAND_166 = {1{`RANDOM}};
  mem_166 = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  mem_167 = _RAND_167[19:0];
  _RAND_168 = {1{`RANDOM}};
  mem_168 = _RAND_168[19:0];
  _RAND_169 = {1{`RANDOM}};
  mem_169 = _RAND_169[19:0];
  _RAND_170 = {1{`RANDOM}};
  mem_170 = _RAND_170[19:0];
  _RAND_171 = {1{`RANDOM}};
  mem_171 = _RAND_171[19:0];
  _RAND_172 = {1{`RANDOM}};
  mem_172 = _RAND_172[19:0];
  _RAND_173 = {1{`RANDOM}};
  mem_173 = _RAND_173[19:0];
  _RAND_174 = {1{`RANDOM}};
  mem_174 = _RAND_174[19:0];
  _RAND_175 = {1{`RANDOM}};
  mem_175 = _RAND_175[19:0];
  _RAND_176 = {1{`RANDOM}};
  mem_176 = _RAND_176[19:0];
  _RAND_177 = {1{`RANDOM}};
  mem_177 = _RAND_177[19:0];
  _RAND_178 = {1{`RANDOM}};
  mem_178 = _RAND_178[19:0];
  _RAND_179 = {1{`RANDOM}};
  mem_179 = _RAND_179[19:0];
  _RAND_180 = {1{`RANDOM}};
  mem_180 = _RAND_180[19:0];
  _RAND_181 = {1{`RANDOM}};
  mem_181 = _RAND_181[19:0];
  _RAND_182 = {1{`RANDOM}};
  mem_182 = _RAND_182[19:0];
  _RAND_183 = {1{`RANDOM}};
  mem_183 = _RAND_183[19:0];
  _RAND_184 = {1{`RANDOM}};
  mem_184 = _RAND_184[19:0];
  _RAND_185 = {1{`RANDOM}};
  mem_185 = _RAND_185[19:0];
  _RAND_186 = {1{`RANDOM}};
  mem_186 = _RAND_186[19:0];
  _RAND_187 = {1{`RANDOM}};
  mem_187 = _RAND_187[19:0];
  _RAND_188 = {1{`RANDOM}};
  mem_188 = _RAND_188[19:0];
  _RAND_189 = {1{`RANDOM}};
  mem_189 = _RAND_189[19:0];
  _RAND_190 = {1{`RANDOM}};
  mem_190 = _RAND_190[19:0];
  _RAND_191 = {1{`RANDOM}};
  mem_191 = _RAND_191[19:0];
  _RAND_192 = {1{`RANDOM}};
  mem_192 = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  mem_193 = _RAND_193[19:0];
  _RAND_194 = {1{`RANDOM}};
  mem_194 = _RAND_194[19:0];
  _RAND_195 = {1{`RANDOM}};
  mem_195 = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  mem_196 = _RAND_196[19:0];
  _RAND_197 = {1{`RANDOM}};
  mem_197 = _RAND_197[19:0];
  _RAND_198 = {1{`RANDOM}};
  mem_198 = _RAND_198[19:0];
  _RAND_199 = {1{`RANDOM}};
  mem_199 = _RAND_199[19:0];
  _RAND_200 = {1{`RANDOM}};
  mem_200 = _RAND_200[19:0];
  _RAND_201 = {1{`RANDOM}};
  mem_201 = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  mem_202 = _RAND_202[19:0];
  _RAND_203 = {1{`RANDOM}};
  mem_203 = _RAND_203[19:0];
  _RAND_204 = {1{`RANDOM}};
  mem_204 = _RAND_204[19:0];
  _RAND_205 = {1{`RANDOM}};
  mem_205 = _RAND_205[19:0];
  _RAND_206 = {1{`RANDOM}};
  mem_206 = _RAND_206[19:0];
  _RAND_207 = {1{`RANDOM}};
  mem_207 = _RAND_207[19:0];
  _RAND_208 = {1{`RANDOM}};
  mem_208 = _RAND_208[19:0];
  _RAND_209 = {1{`RANDOM}};
  mem_209 = _RAND_209[19:0];
  _RAND_210 = {1{`RANDOM}};
  mem_210 = _RAND_210[19:0];
  _RAND_211 = {1{`RANDOM}};
  mem_211 = _RAND_211[19:0];
  _RAND_212 = {1{`RANDOM}};
  mem_212 = _RAND_212[19:0];
  _RAND_213 = {1{`RANDOM}};
  mem_213 = _RAND_213[19:0];
  _RAND_214 = {1{`RANDOM}};
  mem_214 = _RAND_214[19:0];
  _RAND_215 = {1{`RANDOM}};
  mem_215 = _RAND_215[19:0];
  _RAND_216 = {1{`RANDOM}};
  mem_216 = _RAND_216[19:0];
  _RAND_217 = {1{`RANDOM}};
  mem_217 = _RAND_217[19:0];
  _RAND_218 = {1{`RANDOM}};
  mem_218 = _RAND_218[19:0];
  _RAND_219 = {1{`RANDOM}};
  mem_219 = _RAND_219[19:0];
  _RAND_220 = {1{`RANDOM}};
  mem_220 = _RAND_220[19:0];
  _RAND_221 = {1{`RANDOM}};
  mem_221 = _RAND_221[19:0];
  _RAND_222 = {1{`RANDOM}};
  mem_222 = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  mem_223 = _RAND_223[19:0];
  _RAND_224 = {1{`RANDOM}};
  mem_224 = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  mem_225 = _RAND_225[19:0];
  _RAND_226 = {1{`RANDOM}};
  mem_226 = _RAND_226[19:0];
  _RAND_227 = {1{`RANDOM}};
  mem_227 = _RAND_227[19:0];
  _RAND_228 = {1{`RANDOM}};
  mem_228 = _RAND_228[19:0];
  _RAND_229 = {1{`RANDOM}};
  mem_229 = _RAND_229[19:0];
  _RAND_230 = {1{`RANDOM}};
  mem_230 = _RAND_230[19:0];
  _RAND_231 = {1{`RANDOM}};
  mem_231 = _RAND_231[19:0];
  _RAND_232 = {1{`RANDOM}};
  mem_232 = _RAND_232[19:0];
  _RAND_233 = {1{`RANDOM}};
  mem_233 = _RAND_233[19:0];
  _RAND_234 = {1{`RANDOM}};
  mem_234 = _RAND_234[19:0];
  _RAND_235 = {1{`RANDOM}};
  mem_235 = _RAND_235[19:0];
  _RAND_236 = {1{`RANDOM}};
  mem_236 = _RAND_236[19:0];
  _RAND_237 = {1{`RANDOM}};
  mem_237 = _RAND_237[19:0];
  _RAND_238 = {1{`RANDOM}};
  mem_238 = _RAND_238[19:0];
  _RAND_239 = {1{`RANDOM}};
  mem_239 = _RAND_239[19:0];
  _RAND_240 = {1{`RANDOM}};
  mem_240 = _RAND_240[19:0];
  _RAND_241 = {1{`RANDOM}};
  mem_241 = _RAND_241[19:0];
  _RAND_242 = {1{`RANDOM}};
  mem_242 = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  mem_243 = _RAND_243[19:0];
  _RAND_244 = {1{`RANDOM}};
  mem_244 = _RAND_244[19:0];
  _RAND_245 = {1{`RANDOM}};
  mem_245 = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  mem_246 = _RAND_246[19:0];
  _RAND_247 = {1{`RANDOM}};
  mem_247 = _RAND_247[19:0];
  _RAND_248 = {1{`RANDOM}};
  mem_248 = _RAND_248[19:0];
  _RAND_249 = {1{`RANDOM}};
  mem_249 = _RAND_249[19:0];
  _RAND_250 = {1{`RANDOM}};
  mem_250 = _RAND_250[19:0];
  _RAND_251 = {1{`RANDOM}};
  mem_251 = _RAND_251[19:0];
  _RAND_252 = {1{`RANDOM}};
  mem_252 = _RAND_252[19:0];
  _RAND_253 = {1{`RANDOM}};
  mem_253 = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  mem_254 = _RAND_254[19:0];
  _RAND_255 = {1{`RANDOM}};
  mem_255 = _RAND_255[19:0];
  _RAND_256 = {1{`RANDOM}};
  mem_256 = _RAND_256[19:0];
  _RAND_257 = {1{`RANDOM}};
  mem_257 = _RAND_257[19:0];
  _RAND_258 = {1{`RANDOM}};
  mem_258 = _RAND_258[19:0];
  _RAND_259 = {1{`RANDOM}};
  mem_259 = _RAND_259[19:0];
  _RAND_260 = {1{`RANDOM}};
  mem_260 = _RAND_260[19:0];
  _RAND_261 = {1{`RANDOM}};
  mem_261 = _RAND_261[19:0];
  _RAND_262 = {1{`RANDOM}};
  mem_262 = _RAND_262[19:0];
  _RAND_263 = {1{`RANDOM}};
  mem_263 = _RAND_263[19:0];
  _RAND_264 = {1{`RANDOM}};
  mem_264 = _RAND_264[19:0];
  _RAND_265 = {1{`RANDOM}};
  mem_265 = _RAND_265[19:0];
  _RAND_266 = {1{`RANDOM}};
  mem_266 = _RAND_266[19:0];
  _RAND_267 = {1{`RANDOM}};
  mem_267 = _RAND_267[19:0];
  _RAND_268 = {1{`RANDOM}};
  mem_268 = _RAND_268[19:0];
  _RAND_269 = {1{`RANDOM}};
  mem_269 = _RAND_269[19:0];
  _RAND_270 = {1{`RANDOM}};
  mem_270 = _RAND_270[19:0];
  _RAND_271 = {1{`RANDOM}};
  mem_271 = _RAND_271[19:0];
  _RAND_272 = {1{`RANDOM}};
  mem_272 = _RAND_272[19:0];
  _RAND_273 = {1{`RANDOM}};
  mem_273 = _RAND_273[19:0];
  _RAND_274 = {1{`RANDOM}};
  mem_274 = _RAND_274[19:0];
  _RAND_275 = {1{`RANDOM}};
  mem_275 = _RAND_275[19:0];
  _RAND_276 = {1{`RANDOM}};
  mem_276 = _RAND_276[19:0];
  _RAND_277 = {1{`RANDOM}};
  mem_277 = _RAND_277[19:0];
  _RAND_278 = {1{`RANDOM}};
  mem_278 = _RAND_278[19:0];
  _RAND_279 = {1{`RANDOM}};
  mem_279 = _RAND_279[19:0];
  _RAND_280 = {1{`RANDOM}};
  mem_280 = _RAND_280[19:0];
  _RAND_281 = {1{`RANDOM}};
  mem_281 = _RAND_281[19:0];
  _RAND_282 = {1{`RANDOM}};
  mem_282 = _RAND_282[19:0];
  _RAND_283 = {1{`RANDOM}};
  mem_283 = _RAND_283[19:0];
  _RAND_284 = {1{`RANDOM}};
  mem_284 = _RAND_284[19:0];
  _RAND_285 = {1{`RANDOM}};
  mem_285 = _RAND_285[19:0];
  _RAND_286 = {1{`RANDOM}};
  mem_286 = _RAND_286[19:0];
  _RAND_287 = {1{`RANDOM}};
  mem_287 = _RAND_287[19:0];
  _RAND_288 = {1{`RANDOM}};
  mem_288 = _RAND_288[19:0];
  _RAND_289 = {1{`RANDOM}};
  mem_289 = _RAND_289[19:0];
  _RAND_290 = {1{`RANDOM}};
  mem_290 = _RAND_290[19:0];
  _RAND_291 = {1{`RANDOM}};
  mem_291 = _RAND_291[19:0];
  _RAND_292 = {1{`RANDOM}};
  mem_292 = _RAND_292[19:0];
  _RAND_293 = {1{`RANDOM}};
  mem_293 = _RAND_293[19:0];
  _RAND_294 = {1{`RANDOM}};
  mem_294 = _RAND_294[19:0];
  _RAND_295 = {1{`RANDOM}};
  mem_295 = _RAND_295[19:0];
  _RAND_296 = {1{`RANDOM}};
  mem_296 = _RAND_296[19:0];
  _RAND_297 = {1{`RANDOM}};
  mem_297 = _RAND_297[19:0];
  _RAND_298 = {1{`RANDOM}};
  mem_298 = _RAND_298[19:0];
  _RAND_299 = {1{`RANDOM}};
  mem_299 = _RAND_299[19:0];
  _RAND_300 = {1{`RANDOM}};
  mem_300 = _RAND_300[19:0];
  _RAND_301 = {1{`RANDOM}};
  mem_301 = _RAND_301[19:0];
  _RAND_302 = {1{`RANDOM}};
  mem_302 = _RAND_302[19:0];
  _RAND_303 = {1{`RANDOM}};
  mem_303 = _RAND_303[19:0];
  _RAND_304 = {1{`RANDOM}};
  mem_304 = _RAND_304[19:0];
  _RAND_305 = {1{`RANDOM}};
  mem_305 = _RAND_305[19:0];
  _RAND_306 = {1{`RANDOM}};
  mem_306 = _RAND_306[19:0];
  _RAND_307 = {1{`RANDOM}};
  mem_307 = _RAND_307[19:0];
  _RAND_308 = {1{`RANDOM}};
  mem_308 = _RAND_308[19:0];
  _RAND_309 = {1{`RANDOM}};
  mem_309 = _RAND_309[19:0];
  _RAND_310 = {1{`RANDOM}};
  mem_310 = _RAND_310[19:0];
  _RAND_311 = {1{`RANDOM}};
  mem_311 = _RAND_311[19:0];
  _RAND_312 = {1{`RANDOM}};
  mem_312 = _RAND_312[19:0];
  _RAND_313 = {1{`RANDOM}};
  mem_313 = _RAND_313[19:0];
  _RAND_314 = {1{`RANDOM}};
  mem_314 = _RAND_314[19:0];
  _RAND_315 = {1{`RANDOM}};
  mem_315 = _RAND_315[19:0];
  _RAND_316 = {1{`RANDOM}};
  mem_316 = _RAND_316[19:0];
  _RAND_317 = {1{`RANDOM}};
  mem_317 = _RAND_317[19:0];
  _RAND_318 = {1{`RANDOM}};
  mem_318 = _RAND_318[19:0];
  _RAND_319 = {1{`RANDOM}};
  mem_319 = _RAND_319[19:0];
  _RAND_320 = {1{`RANDOM}};
  mem_320 = _RAND_320[19:0];
  _RAND_321 = {1{`RANDOM}};
  mem_321 = _RAND_321[19:0];
  _RAND_322 = {1{`RANDOM}};
  mem_322 = _RAND_322[19:0];
  _RAND_323 = {1{`RANDOM}};
  mem_323 = _RAND_323[19:0];
  _RAND_324 = {1{`RANDOM}};
  mem_324 = _RAND_324[19:0];
  _RAND_325 = {1{`RANDOM}};
  mem_325 = _RAND_325[19:0];
  _RAND_326 = {1{`RANDOM}};
  mem_326 = _RAND_326[19:0];
  _RAND_327 = {1{`RANDOM}};
  mem_327 = _RAND_327[19:0];
  _RAND_328 = {1{`RANDOM}};
  mem_328 = _RAND_328[19:0];
  _RAND_329 = {1{`RANDOM}};
  mem_329 = _RAND_329[19:0];
  _RAND_330 = {1{`RANDOM}};
  mem_330 = _RAND_330[19:0];
  _RAND_331 = {1{`RANDOM}};
  mem_331 = _RAND_331[19:0];
  _RAND_332 = {1{`RANDOM}};
  mem_332 = _RAND_332[19:0];
  _RAND_333 = {1{`RANDOM}};
  mem_333 = _RAND_333[19:0];
  _RAND_334 = {1{`RANDOM}};
  mem_334 = _RAND_334[19:0];
  _RAND_335 = {1{`RANDOM}};
  mem_335 = _RAND_335[19:0];
  _RAND_336 = {1{`RANDOM}};
  mem_336 = _RAND_336[19:0];
  _RAND_337 = {1{`RANDOM}};
  mem_337 = _RAND_337[19:0];
  _RAND_338 = {1{`RANDOM}};
  mem_338 = _RAND_338[19:0];
  _RAND_339 = {1{`RANDOM}};
  mem_339 = _RAND_339[19:0];
  _RAND_340 = {1{`RANDOM}};
  mem_340 = _RAND_340[19:0];
  _RAND_341 = {1{`RANDOM}};
  mem_341 = _RAND_341[19:0];
  _RAND_342 = {1{`RANDOM}};
  mem_342 = _RAND_342[19:0];
  _RAND_343 = {1{`RANDOM}};
  mem_343 = _RAND_343[19:0];
  _RAND_344 = {1{`RANDOM}};
  mem_344 = _RAND_344[19:0];
  _RAND_345 = {1{`RANDOM}};
  mem_345 = _RAND_345[19:0];
  _RAND_346 = {1{`RANDOM}};
  mem_346 = _RAND_346[19:0];
  _RAND_347 = {1{`RANDOM}};
  mem_347 = _RAND_347[19:0];
  _RAND_348 = {1{`RANDOM}};
  mem_348 = _RAND_348[19:0];
  _RAND_349 = {1{`RANDOM}};
  mem_349 = _RAND_349[19:0];
  _RAND_350 = {1{`RANDOM}};
  mem_350 = _RAND_350[19:0];
  _RAND_351 = {1{`RANDOM}};
  mem_351 = _RAND_351[19:0];
  _RAND_352 = {1{`RANDOM}};
  mem_352 = _RAND_352[19:0];
  _RAND_353 = {1{`RANDOM}};
  mem_353 = _RAND_353[19:0];
  _RAND_354 = {1{`RANDOM}};
  mem_354 = _RAND_354[19:0];
  _RAND_355 = {1{`RANDOM}};
  mem_355 = _RAND_355[19:0];
  _RAND_356 = {1{`RANDOM}};
  mem_356 = _RAND_356[19:0];
  _RAND_357 = {1{`RANDOM}};
  mem_357 = _RAND_357[19:0];
  _RAND_358 = {1{`RANDOM}};
  mem_358 = _RAND_358[19:0];
  _RAND_359 = {1{`RANDOM}};
  mem_359 = _RAND_359[19:0];
  _RAND_360 = {1{`RANDOM}};
  mem_360 = _RAND_360[19:0];
  _RAND_361 = {1{`RANDOM}};
  mem_361 = _RAND_361[19:0];
  _RAND_362 = {1{`RANDOM}};
  mem_362 = _RAND_362[19:0];
  _RAND_363 = {1{`RANDOM}};
  mem_363 = _RAND_363[19:0];
  _RAND_364 = {1{`RANDOM}};
  mem_364 = _RAND_364[19:0];
  _RAND_365 = {1{`RANDOM}};
  mem_365 = _RAND_365[19:0];
  _RAND_366 = {1{`RANDOM}};
  mem_366 = _RAND_366[19:0];
  _RAND_367 = {1{`RANDOM}};
  mem_367 = _RAND_367[19:0];
  _RAND_368 = {1{`RANDOM}};
  mem_368 = _RAND_368[19:0];
  _RAND_369 = {1{`RANDOM}};
  mem_369 = _RAND_369[19:0];
  _RAND_370 = {1{`RANDOM}};
  mem_370 = _RAND_370[19:0];
  _RAND_371 = {1{`RANDOM}};
  mem_371 = _RAND_371[19:0];
  _RAND_372 = {1{`RANDOM}};
  mem_372 = _RAND_372[19:0];
  _RAND_373 = {1{`RANDOM}};
  mem_373 = _RAND_373[19:0];
  _RAND_374 = {1{`RANDOM}};
  mem_374 = _RAND_374[19:0];
  _RAND_375 = {1{`RANDOM}};
  mem_375 = _RAND_375[19:0];
  _RAND_376 = {1{`RANDOM}};
  mem_376 = _RAND_376[19:0];
  _RAND_377 = {1{`RANDOM}};
  mem_377 = _RAND_377[19:0];
  _RAND_378 = {1{`RANDOM}};
  mem_378 = _RAND_378[19:0];
  _RAND_379 = {1{`RANDOM}};
  mem_379 = _RAND_379[19:0];
  _RAND_380 = {1{`RANDOM}};
  mem_380 = _RAND_380[19:0];
  _RAND_381 = {1{`RANDOM}};
  mem_381 = _RAND_381[19:0];
  _RAND_382 = {1{`RANDOM}};
  mem_382 = _RAND_382[19:0];
  _RAND_383 = {1{`RANDOM}};
  mem_383 = _RAND_383[19:0];
  _RAND_384 = {1{`RANDOM}};
  mem_384 = _RAND_384[19:0];
  _RAND_385 = {1{`RANDOM}};
  mem_385 = _RAND_385[19:0];
  _RAND_386 = {1{`RANDOM}};
  mem_386 = _RAND_386[19:0];
  _RAND_387 = {1{`RANDOM}};
  mem_387 = _RAND_387[19:0];
  _RAND_388 = {1{`RANDOM}};
  mem_388 = _RAND_388[19:0];
  _RAND_389 = {1{`RANDOM}};
  mem_389 = _RAND_389[19:0];
  _RAND_390 = {1{`RANDOM}};
  mem_390 = _RAND_390[19:0];
  _RAND_391 = {1{`RANDOM}};
  mem_391 = _RAND_391[19:0];
  _RAND_392 = {1{`RANDOM}};
  mem_392 = _RAND_392[19:0];
  _RAND_393 = {1{`RANDOM}};
  mem_393 = _RAND_393[19:0];
  _RAND_394 = {1{`RANDOM}};
  mem_394 = _RAND_394[19:0];
  _RAND_395 = {1{`RANDOM}};
  mem_395 = _RAND_395[19:0];
  _RAND_396 = {1{`RANDOM}};
  mem_396 = _RAND_396[19:0];
  _RAND_397 = {1{`RANDOM}};
  mem_397 = _RAND_397[19:0];
  _RAND_398 = {1{`RANDOM}};
  mem_398 = _RAND_398[19:0];
  _RAND_399 = {1{`RANDOM}};
  mem_399 = _RAND_399[19:0];
  _RAND_400 = {1{`RANDOM}};
  mem_400 = _RAND_400[19:0];
  _RAND_401 = {1{`RANDOM}};
  mem_401 = _RAND_401[19:0];
  _RAND_402 = {1{`RANDOM}};
  mem_402 = _RAND_402[19:0];
  _RAND_403 = {1{`RANDOM}};
  mem_403 = _RAND_403[19:0];
  _RAND_404 = {1{`RANDOM}};
  mem_404 = _RAND_404[19:0];
  _RAND_405 = {1{`RANDOM}};
  mem_405 = _RAND_405[19:0];
  _RAND_406 = {1{`RANDOM}};
  mem_406 = _RAND_406[19:0];
  _RAND_407 = {1{`RANDOM}};
  mem_407 = _RAND_407[19:0];
  _RAND_408 = {1{`RANDOM}};
  mem_408 = _RAND_408[19:0];
  _RAND_409 = {1{`RANDOM}};
  mem_409 = _RAND_409[19:0];
  _RAND_410 = {1{`RANDOM}};
  mem_410 = _RAND_410[19:0];
  _RAND_411 = {1{`RANDOM}};
  mem_411 = _RAND_411[19:0];
  _RAND_412 = {1{`RANDOM}};
  mem_412 = _RAND_412[19:0];
  _RAND_413 = {1{`RANDOM}};
  mem_413 = _RAND_413[19:0];
  _RAND_414 = {1{`RANDOM}};
  mem_414 = _RAND_414[19:0];
  _RAND_415 = {1{`RANDOM}};
  mem_415 = _RAND_415[19:0];
  _RAND_416 = {1{`RANDOM}};
  mem_416 = _RAND_416[19:0];
  _RAND_417 = {1{`RANDOM}};
  mem_417 = _RAND_417[19:0];
  _RAND_418 = {1{`RANDOM}};
  mem_418 = _RAND_418[19:0];
  _RAND_419 = {1{`RANDOM}};
  mem_419 = _RAND_419[19:0];
  _RAND_420 = {1{`RANDOM}};
  mem_420 = _RAND_420[19:0];
  _RAND_421 = {1{`RANDOM}};
  mem_421 = _RAND_421[19:0];
  _RAND_422 = {1{`RANDOM}};
  mem_422 = _RAND_422[19:0];
  _RAND_423 = {1{`RANDOM}};
  mem_423 = _RAND_423[19:0];
  _RAND_424 = {1{`RANDOM}};
  mem_424 = _RAND_424[19:0];
  _RAND_425 = {1{`RANDOM}};
  mem_425 = _RAND_425[19:0];
  _RAND_426 = {1{`RANDOM}};
  mem_426 = _RAND_426[19:0];
  _RAND_427 = {1{`RANDOM}};
  mem_427 = _RAND_427[19:0];
  _RAND_428 = {1{`RANDOM}};
  mem_428 = _RAND_428[19:0];
  _RAND_429 = {1{`RANDOM}};
  mem_429 = _RAND_429[19:0];
  _RAND_430 = {1{`RANDOM}};
  mem_430 = _RAND_430[19:0];
  _RAND_431 = {1{`RANDOM}};
  mem_431 = _RAND_431[19:0];
  _RAND_432 = {1{`RANDOM}};
  mem_432 = _RAND_432[19:0];
  _RAND_433 = {1{`RANDOM}};
  mem_433 = _RAND_433[19:0];
  _RAND_434 = {1{`RANDOM}};
  mem_434 = _RAND_434[19:0];
  _RAND_435 = {1{`RANDOM}};
  mem_435 = _RAND_435[19:0];
  _RAND_436 = {1{`RANDOM}};
  mem_436 = _RAND_436[19:0];
  _RAND_437 = {1{`RANDOM}};
  mem_437 = _RAND_437[19:0];
  _RAND_438 = {1{`RANDOM}};
  mem_438 = _RAND_438[19:0];
  _RAND_439 = {1{`RANDOM}};
  mem_439 = _RAND_439[19:0];
  _RAND_440 = {1{`RANDOM}};
  mem_440 = _RAND_440[19:0];
  _RAND_441 = {1{`RANDOM}};
  mem_441 = _RAND_441[19:0];
  _RAND_442 = {1{`RANDOM}};
  mem_442 = _RAND_442[19:0];
  _RAND_443 = {1{`RANDOM}};
  mem_443 = _RAND_443[19:0];
  _RAND_444 = {1{`RANDOM}};
  mem_444 = _RAND_444[19:0];
  _RAND_445 = {1{`RANDOM}};
  mem_445 = _RAND_445[19:0];
  _RAND_446 = {1{`RANDOM}};
  mem_446 = _RAND_446[19:0];
  _RAND_447 = {1{`RANDOM}};
  mem_447 = _RAND_447[19:0];
  _RAND_448 = {1{`RANDOM}};
  mem_448 = _RAND_448[19:0];
  _RAND_449 = {1{`RANDOM}};
  mem_449 = _RAND_449[19:0];
  _RAND_450 = {1{`RANDOM}};
  mem_450 = _RAND_450[19:0];
  _RAND_451 = {1{`RANDOM}};
  mem_451 = _RAND_451[19:0];
  _RAND_452 = {1{`RANDOM}};
  mem_452 = _RAND_452[19:0];
  _RAND_453 = {1{`RANDOM}};
  mem_453 = _RAND_453[19:0];
  _RAND_454 = {1{`RANDOM}};
  mem_454 = _RAND_454[19:0];
  _RAND_455 = {1{`RANDOM}};
  mem_455 = _RAND_455[19:0];
  _RAND_456 = {1{`RANDOM}};
  mem_456 = _RAND_456[19:0];
  _RAND_457 = {1{`RANDOM}};
  mem_457 = _RAND_457[19:0];
  _RAND_458 = {1{`RANDOM}};
  mem_458 = _RAND_458[19:0];
  _RAND_459 = {1{`RANDOM}};
  mem_459 = _RAND_459[19:0];
  _RAND_460 = {1{`RANDOM}};
  mem_460 = _RAND_460[19:0];
  _RAND_461 = {1{`RANDOM}};
  mem_461 = _RAND_461[19:0];
  _RAND_462 = {1{`RANDOM}};
  mem_462 = _RAND_462[19:0];
  _RAND_463 = {1{`RANDOM}};
  mem_463 = _RAND_463[19:0];
  _RAND_464 = {1{`RANDOM}};
  mem_464 = _RAND_464[19:0];
  _RAND_465 = {1{`RANDOM}};
  mem_465 = _RAND_465[19:0];
  _RAND_466 = {1{`RANDOM}};
  mem_466 = _RAND_466[19:0];
  _RAND_467 = {1{`RANDOM}};
  mem_467 = _RAND_467[19:0];
  _RAND_468 = {1{`RANDOM}};
  mem_468 = _RAND_468[19:0];
  _RAND_469 = {1{`RANDOM}};
  mem_469 = _RAND_469[19:0];
  _RAND_470 = {1{`RANDOM}};
  mem_470 = _RAND_470[19:0];
  _RAND_471 = {1{`RANDOM}};
  mem_471 = _RAND_471[19:0];
  _RAND_472 = {1{`RANDOM}};
  mem_472 = _RAND_472[19:0];
  _RAND_473 = {1{`RANDOM}};
  mem_473 = _RAND_473[19:0];
  _RAND_474 = {1{`RANDOM}};
  mem_474 = _RAND_474[19:0];
  _RAND_475 = {1{`RANDOM}};
  mem_475 = _RAND_475[19:0];
  _RAND_476 = {1{`RANDOM}};
  mem_476 = _RAND_476[19:0];
  _RAND_477 = {1{`RANDOM}};
  mem_477 = _RAND_477[19:0];
  _RAND_478 = {1{`RANDOM}};
  mem_478 = _RAND_478[19:0];
  _RAND_479 = {1{`RANDOM}};
  mem_479 = _RAND_479[19:0];
  _RAND_480 = {1{`RANDOM}};
  mem_480 = _RAND_480[19:0];
  _RAND_481 = {1{`RANDOM}};
  mem_481 = _RAND_481[19:0];
  _RAND_482 = {1{`RANDOM}};
  mem_482 = _RAND_482[19:0];
  _RAND_483 = {1{`RANDOM}};
  mem_483 = _RAND_483[19:0];
  _RAND_484 = {1{`RANDOM}};
  mem_484 = _RAND_484[19:0];
  _RAND_485 = {1{`RANDOM}};
  mem_485 = _RAND_485[19:0];
  _RAND_486 = {1{`RANDOM}};
  mem_486 = _RAND_486[19:0];
  _RAND_487 = {1{`RANDOM}};
  mem_487 = _RAND_487[19:0];
  _RAND_488 = {1{`RANDOM}};
  mem_488 = _RAND_488[19:0];
  _RAND_489 = {1{`RANDOM}};
  mem_489 = _RAND_489[19:0];
  _RAND_490 = {1{`RANDOM}};
  mem_490 = _RAND_490[19:0];
  _RAND_491 = {1{`RANDOM}};
  mem_491 = _RAND_491[19:0];
  _RAND_492 = {1{`RANDOM}};
  mem_492 = _RAND_492[19:0];
  _RAND_493 = {1{`RANDOM}};
  mem_493 = _RAND_493[19:0];
  _RAND_494 = {1{`RANDOM}};
  mem_494 = _RAND_494[19:0];
  _RAND_495 = {1{`RANDOM}};
  mem_495 = _RAND_495[19:0];
  _RAND_496 = {1{`RANDOM}};
  mem_496 = _RAND_496[19:0];
  _RAND_497 = {1{`RANDOM}};
  mem_497 = _RAND_497[19:0];
  _RAND_498 = {1{`RANDOM}};
  mem_498 = _RAND_498[19:0];
  _RAND_499 = {1{`RANDOM}};
  mem_499 = _RAND_499[19:0];
  _RAND_500 = {1{`RANDOM}};
  mem_500 = _RAND_500[19:0];
  _RAND_501 = {1{`RANDOM}};
  mem_501 = _RAND_501[19:0];
  _RAND_502 = {1{`RANDOM}};
  mem_502 = _RAND_502[19:0];
  _RAND_503 = {1{`RANDOM}};
  mem_503 = _RAND_503[19:0];
  _RAND_504 = {1{`RANDOM}};
  mem_504 = _RAND_504[19:0];
  _RAND_505 = {1{`RANDOM}};
  mem_505 = _RAND_505[19:0];
  _RAND_506 = {1{`RANDOM}};
  mem_506 = _RAND_506[19:0];
  _RAND_507 = {1{`RANDOM}};
  mem_507 = _RAND_507[19:0];
  _RAND_508 = {1{`RANDOM}};
  mem_508 = _RAND_508[19:0];
  _RAND_509 = {1{`RANDOM}};
  mem_509 = _RAND_509[19:0];
  _RAND_510 = {1{`RANDOM}};
  mem_510 = _RAND_510[19:0];
  _RAND_511 = {1{`RANDOM}};
  mem_511 = _RAND_511[19:0];
  _RAND_512 = {1{`RANDOM}};
  io_douta_REG = _RAND_512[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM_3(
  input         clock,
  input         reset,
  input         io_web,
  input  [8:0]  io_addra,
  input  [8:0]  io_addrb,
  input  [19:0] io_dinb,
  output [19:0] io_douta
);
  wire  sim_dual_port_bram_clock; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_reset; // @[RAMWrapper.scala 30:36]
  wire  sim_dual_port_bram_io_web; // @[RAMWrapper.scala 30:36]
  wire [8:0] sim_dual_port_bram_io_addra; // @[RAMWrapper.scala 30:36]
  wire [8:0] sim_dual_port_bram_io_addrb; // @[RAMWrapper.scala 30:36]
  wire [19:0] sim_dual_port_bram_io_dinb; // @[RAMWrapper.scala 30:36]
  wire [19:0] sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 30:36]
  SimDualPortBRAM_3 sim_dual_port_bram ( // @[RAMWrapper.scala 30:36]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_web(sim_dual_port_bram_io_web),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dinb(sim_dual_port_bram_io_dinb),
    .io_douta(sim_dual_port_bram_io_douta)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_web = io_web; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAMWrapper.scala 31:27]
  assign sim_dual_port_bram_io_dinb = io_dinb; // @[RAMWrapper.scala 31:27]
endmodule
module MetaDataBRAM(
  input         clock,
  input         reset,
  input  [8:0]  io_index_fetch,
  input  [8:0]  io_index_update,
  input  [17:0] io_tag_update,
  input         io_update,
  input         io_write,
  output        io_hit,
  output [17:0] io_tag_fetch,
  output        io_dirty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  blk_clock; // @[Dcache.scala 27:19]
  wire  blk_reset; // @[Dcache.scala 27:19]
  wire  blk_io_web; // @[Dcache.scala 27:19]
  wire [8:0] blk_io_addra; // @[Dcache.scala 27:19]
  wire [8:0] blk_io_addrb; // @[Dcache.scala 27:19]
  wire [19:0] blk_io_dinb; // @[Dcache.scala 27:19]
  wire [19:0] blk_io_douta; // @[Dcache.scala 27:19]
  reg  dout_REG; // @[Dcache.scala 30:25]
  reg [19:0] dout_REG_1; // @[Dcache.scala 30:79]
  wire [19:0] dout = dout_REG ? dout_REG_1 : blk_io_douta; // @[Dcache.scala 30:17]
  wire  v = dout[18]; // @[Dcache.scala 31:15]
  wire [17:0] tag = dout[17:0]; // @[Dcache.scala 32:17]
  wire [1:0] blk_io_dinb_hi = {io_write,1'h1}; // @[Cat.scala 30:58]
  DualPortBRAM_3 blk ( // @[Dcache.scala 27:19]
    .clock(blk_clock),
    .reset(blk_reset),
    .io_web(blk_io_web),
    .io_addra(blk_io_addra),
    .io_addrb(blk_io_addrb),
    .io_dinb(blk_io_dinb),
    .io_douta(blk_io_douta)
  );
  assign io_hit = v & io_tag_update == tag; // @[Dcache.scala 51:21]
  assign io_tag_fetch = dout[17:0]; // @[Dcache.scala 32:17]
  assign io_dirty = dout[19]; // @[Dcache.scala 50:23]
  assign blk_clock = clock;
  assign blk_reset = reset;
  assign blk_io_web = io_update; // @[Dcache.scala 46:16]
  assign blk_io_addra = io_index_fetch; // @[Dcache.scala 42:16]
  assign blk_io_addrb = io_index_update; // @[Dcache.scala 47:16]
  assign blk_io_dinb = {blk_io_dinb_hi,io_tag_update}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    dout_REG <= blk_io_web & blk_io_addra == blk_io_addrb; // @[Dcache.scala 30:37]
    dout_REG_1 <= blk_io_dinb; // @[Dcache.scala 30:79]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dout_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dout_REG_1 = _RAND_1[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DcacheDP(
  input          clock,
  input          reset,
  input          io_cpu_req_valid,
  input  [31:0]  io_cpu_req_bits_addr,
  input  [63:0]  io_cpu_req_bits_wdata,
  input          io_cpu_req_bits_wen,
  input  [2:0]   io_cpu_req_bits_mtype,
  output         io_cpu_resp_valid,
  output [31:0]  io_cpu_resp_bits_rdata_0,
  output [31:0]  io_cpu_resp_bits_rdata_1,
  output         io_bar_req_valid,
  output         io_bar_req_wen,
  output [31:0]  io_bar_req_addr,
  output [255:0] io_bar_req_data,
  output [2:0]   io_bar_req_mtype,
  input          io_bar_resp_valid,
  input  [255:0] io_bar_resp_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  data_clock; // @[Dcache.scala 66:20]
  wire  data_reset; // @[Dcache.scala 66:20]
  wire  data_io_web; // @[Dcache.scala 66:20]
  wire [8:0] data_io_addra; // @[Dcache.scala 66:20]
  wire [8:0] data_io_addrb; // @[Dcache.scala 66:20]
  wire [255:0] data_io_dinb; // @[Dcache.scala 66:20]
  wire [255:0] data_io_douta; // @[Dcache.scala 66:20]
  wire  meta_clock; // @[Dcache.scala 67:20]
  wire  meta_reset; // @[Dcache.scala 67:20]
  wire [8:0] meta_io_index_fetch; // @[Dcache.scala 67:20]
  wire [8:0] meta_io_index_update; // @[Dcache.scala 67:20]
  wire [17:0] meta_io_tag_update; // @[Dcache.scala 67:20]
  wire  meta_io_update; // @[Dcache.scala 67:20]
  wire  meta_io_write; // @[Dcache.scala 67:20]
  wire  meta_io_hit; // @[Dcache.scala 67:20]
  wire [17:0] meta_io_tag_fetch; // @[Dcache.scala 67:20]
  wire  meta_io_dirty; // @[Dcache.scala 67:20]
  wire [8:0] df_index = io_cpu_req_bits_addr[13:5]; // @[Dcache.scala 74:49]
  wire [17:0] df_tag = io_cpu_req_bits_addr[31:14]; // @[Dcache.scala 75:49]
  wire [1:0] df_offset = io_cpu_req_bits_addr[4:3]; // @[Dcache.scala 76:49]
  reg  wb_valid; // @[Dcache.scala 97:31]
  reg  wb_state; // @[Dcache.scala 201:25]
  wire  _T_22 = ~wb_state; // @[Conditional.scala 37:30]
  wire  wb_write_cache = wb_valid & wb_state & io_bar_resp_valid; // @[Dcache.scala 203:58]
  wire  _GEN_53 = wb_state & wb_write_cache; // @[Conditional.scala 39:67 Dcache.scala 244:23 Dcache.scala 236:17]
  wire  _GEN_56 = _T_22 ? 1'h0 : _GEN_53; // @[Conditional.scala 40:58 Dcache.scala 236:17]
  wire  wb_resp_valid = wb_valid & _GEN_56; // @[Dcache.scala 237:19 Dcache.scala 236:17]
  wire  wb_stall = wb_valid & ~wb_resp_valid; // @[Dcache.scala 105:33]
  wire  _dp_index_T = ~wb_stall; // @[Dcache.scala 83:49]
  reg [8:0] dp_index; // @[Reg.scala 15:16]
  reg [17:0] dp_tag; // @[Reg.scala 15:16]
  reg [1:0] dp_offset; // @[Reg.scala 15:16]
  reg [31:0] dp_req_addr; // @[Reg.scala 15:16]
  reg [63:0] dp_req_wdata; // @[Reg.scala 15:16]
  reg  dp_req_wen; // @[Reg.scala 15:16]
  reg [2:0] dp_req_mtype; // @[Reg.scala 15:16]
  reg  dp_valid; // @[Dcache.scala 87:36]
  wire  dp_resp_valid = dp_valid & meta_io_hit; // @[Dcache.scala 88:38]
  reg  dp_mmio_valid; // @[Reg.scala 15:16]
  wire  _dp_mmio_stall_T = ~io_bar_resp_valid; // @[Dcache.scala 128:37]
  wire  dp_mmio_stall = dp_mmio_valid & ~io_bar_resp_valid; // @[Dcache.scala 128:34]
  wire  _dp_mmio_valid_T = ~dp_mmio_stall; // @[Dcache.scala 90:54]
  wire  df_mmio_valid = (dp_resp_valid | ~dp_valid & ~wb_valid) & ~io_cpu_req_bits_addr[31] & io_cpu_req_valid; // @[Dcache.scala 133:101]
  reg [31:0] dp_mmio_req_addr; // @[Reg.scala 15:16]
  reg [63:0] dp_mmio_req_wdata; // @[Reg.scala 15:16]
  reg  dp_mmio_req_wen; // @[Reg.scala 15:16]
  reg [2:0] dp_mmio_req_mtype; // @[Reg.scala 15:16]
  reg [255:0] wb_dirty_data; // @[Dcache.scala 95:27]
  reg [31:0] wb_dirty_addr; // @[Dcache.scala 96:27]
  reg [63:0] wb_req_wdata; // @[Dcache.scala 99:31]
  reg  wb_req_wen; // @[Dcache.scala 99:31]
  reg [8:0] wb_index; // @[Dcache.scala 100:27]
  reg [17:0] wb_tag; // @[Dcache.scala 101:27]
  reg [4:0] wb_offset; // @[Dcache.scala 102:27]
  wire [31:0] wb_refill_addr = {wb_tag,wb_index,5'h0}; // @[Cat.scala 30:58]
  reg [63:0] wb_mask; // @[Dcache.scala 109:27]
  reg [5:0] wb_shift; // @[Dcache.scala 110:27]
  wire  dp_mmio_resp_valid = dp_mmio_valid & io_bar_resp_valid; // @[Dcache.scala 137:39]
  reg  REG; // @[Dcache.scala 153:31]
  wire [255:0] _WIRE_1 = data_io_dinb;
  reg [63:0] REG_1_0; // @[Dcache.scala 154:12]
  reg [63:0] REG_1_1; // @[Dcache.scala 154:12]
  reg [63:0] REG_1_2; // @[Dcache.scala 154:12]
  reg [63:0] REG_1_3; // @[Dcache.scala 154:12]
  wire [255:0] _WIRE_3 = data_io_douta;
  wire [63:0] dp_fetch_line_0 = REG ? REG_1_0 : _WIRE_3[63:0]; // @[Dcache.scala 153:23]
  wire [63:0] dp_fetch_line_1 = REG ? REG_1_1 : _WIRE_3[127:64]; // @[Dcache.scala 153:23]
  wire [63:0] dp_fetch_line_2 = REG ? REG_1_2 : _WIRE_3[191:128]; // @[Dcache.scala 153:23]
  wire [63:0] dp_fetch_line_3 = REG ? REG_1_3 : _WIRE_3[255:192]; // @[Dcache.scala 153:23]
  wire  _dp_valid_T_1 = dp_valid & ~meta_io_hit; // @[Dcache.scala 157:33]
  wire [63:0] _dp_mask_T_1 = 3'h1 == dp_req_mtype ? 64'hffff : 64'hffffffffffffffff; // @[Mux.scala 80:57]
  wire [63:0] _dp_mask_T_3 = 3'h0 == dp_req_mtype ? 64'hff : _dp_mask_T_1; // @[Mux.scala 80:57]
  wire [63:0] dp_mask = 3'h2 == dp_req_mtype ? 64'hffffffff : _dp_mask_T_3; // @[Mux.scala 80:57]
  wire [5:0] dp_shift = {dp_req_addr[2:0], 3'h0}; // @[Dcache.scala 172:51]
  wire [63:0] _dp_write_word_T = dp_mask & dp_req_wdata; // @[Dcache.scala 173:33]
  wire [126:0] _GEN_60 = {{63'd0}, _dp_write_word_T}; // @[Dcache.scala 173:49]
  wire [126:0] _dp_write_word_T_1 = _GEN_60 << dp_shift; // @[Dcache.scala 173:49]
  wire [126:0] _GEN_61 = {{63'd0}, dp_mask}; // @[Dcache.scala 173:85]
  wire [126:0] _dp_write_word_T_2 = _GEN_61 << dp_shift; // @[Dcache.scala 173:85]
  wire [126:0] _dp_write_word_T_3 = ~_dp_write_word_T_2; // @[Dcache.scala 173:75]
  wire [63:0] _GEN_17 = 2'h1 == dp_offset ? dp_fetch_line_1 : dp_fetch_line_0; // @[Dcache.scala 173:108 Dcache.scala 173:108]
  wire [63:0] _GEN_18 = 2'h2 == dp_offset ? dp_fetch_line_2 : _GEN_17; // @[Dcache.scala 173:108 Dcache.scala 173:108]
  wire [63:0] _GEN_19 = 2'h3 == dp_offset ? dp_fetch_line_3 : _GEN_18; // @[Dcache.scala 173:108 Dcache.scala 173:108]
  wire [126:0] _GEN_62 = {{63'd0}, _GEN_19}; // @[Dcache.scala 173:108]
  wire [126:0] _dp_write_word_T_4 = _dp_write_word_T_3 & _GEN_62; // @[Dcache.scala 173:108]
  wire [126:0] dp_write_word = _dp_write_word_T_1 | _dp_write_word_T_4; // @[Dcache.scala 173:71]
  wire [31:0] UNCACHED_RESP_RDATA_hi = io_bar_resp_data[31:0]; // @[Dcache.scala 174:67]
  wire [63:0] UNCACHED_RESP_RDATA = {UNCACHED_RESP_RDATA_hi,UNCACHED_RESP_RDATA_hi}; // @[Cat.scala 30:58]
  wire [63:0] dp_write_line_0 = 2'h0 == dp_offset ? dp_write_word[63:0] : dp_fetch_line_0; // @[Dcache.scala 176:28 Dcache.scala 176:28 Dcache.scala 175:17]
  wire [63:0] dp_write_line_1 = 2'h1 == dp_offset ? dp_write_word[63:0] : dp_fetch_line_1; // @[Dcache.scala 176:28 Dcache.scala 176:28 Dcache.scala 175:17]
  wire [63:0] dp_write_line_2 = 2'h2 == dp_offset ? dp_write_word[63:0] : dp_fetch_line_2; // @[Dcache.scala 176:28 Dcache.scala 176:28 Dcache.scala 175:17]
  wire [63:0] dp_write_line_3 = 2'h3 == dp_offset ? dp_write_word[63:0] : dp_fetch_line_3; // @[Dcache.scala 176:28 Dcache.scala 176:28 Dcache.scala 175:17]
  wire [63:0] _T_12 = dp_mmio_valid ? UNCACHED_RESP_RDATA : _GEN_19; // @[Dcache.scala 183:8]
  wire [63:0] wb_refill_line_0 = io_bar_resp_data[63:0]; // @[Dcache.scala 215:48]
  wire [63:0] wb_refill_line_1 = io_bar_resp_data[127:64]; // @[Dcache.scala 215:48]
  wire [63:0] _GEN_25 = 2'h1 == wb_offset[1:0] ? wb_refill_line_1 : wb_refill_line_0; // @[Dcache.scala 182:35 Dcache.scala 182:35]
  wire [63:0] wb_refill_line_2 = io_bar_resp_data[191:128]; // @[Dcache.scala 215:48]
  wire [63:0] _GEN_26 = 2'h2 == wb_offset[1:0] ? wb_refill_line_2 : _GEN_25; // @[Dcache.scala 182:35 Dcache.scala 182:35]
  wire [63:0] wb_refill_line_3 = io_bar_resp_data[255:192]; // @[Dcache.scala 215:48]
  wire [63:0] _GEN_27 = 2'h3 == wb_offset[1:0] ? wb_refill_line_3 : _GEN_26; // @[Dcache.scala 182:35 Dcache.scala 182:35]
  wire [63:0] _T_13 = wb_valid ? _GEN_27 : _T_12; // @[Dcache.scala 182:35]
  wire  _data_io_web_T_1 = dp_resp_valid & dp_req_wen; // @[Dcache.scala 186:74]
  wire [63:0] _wb_write_word_T = wb_mask & wb_req_wdata; // @[Dcache.scala 233:33]
  wire [126:0] _GEN_63 = {{63'd0}, _wb_write_word_T}; // @[Dcache.scala 233:49]
  wire [126:0] _wb_write_word_T_1 = _GEN_63 << wb_shift; // @[Dcache.scala 233:49]
  wire [126:0] _GEN_64 = {{63'd0}, wb_mask}; // @[Dcache.scala 233:85]
  wire [126:0] _wb_write_word_T_2 = _GEN_64 << wb_shift; // @[Dcache.scala 233:85]
  wire [126:0] _wb_write_word_T_3 = ~_wb_write_word_T_2; // @[Dcache.scala 233:75]
  wire [126:0] _GEN_65 = {{63'd0}, _GEN_27}; // @[Dcache.scala 233:108]
  wire [126:0] _wb_write_word_T_5 = _wb_write_word_T_3 & _GEN_65; // @[Dcache.scala 233:108]
  wire [126:0] wb_write_word = _wb_write_word_T_1 | _wb_write_word_T_5; // @[Dcache.scala 233:71]
  wire [63:0] wb_write_line_1 = 2'h1 == wb_offset[1:0] ? wb_write_word[63:0] : wb_refill_line_1; // @[Dcache.scala 235:28 Dcache.scala 235:28 Dcache.scala 234:17]
  wire [63:0] wb_write_line_0 = 2'h0 == wb_offset[1:0] ? wb_write_word[63:0] : wb_refill_line_0; // @[Dcache.scala 235:28 Dcache.scala 235:28 Dcache.scala 234:17]
  wire [63:0] wb_write_line_3 = 2'h3 == wb_offset[1:0] ? wb_write_word[63:0] : wb_refill_line_3; // @[Dcache.scala 235:28 Dcache.scala 235:28 Dcache.scala 234:17]
  wire [63:0] wb_write_line_2 = 2'h2 == wb_offset[1:0] ? wb_write_word[63:0] : wb_refill_line_2; // @[Dcache.scala 235:28 Dcache.scala 235:28 Dcache.scala 234:17]
  wire [255:0] _data_io_dinb_T = {wb_write_line_3,wb_write_line_2,wb_write_line_1,wb_write_line_0}; // @[Dcache.scala 187:70]
  wire [255:0] _data_io_dinb_T_1 = wb_req_wen ? _data_io_dinb_T : io_bar_resp_data; // @[Dcache.scala 187:37]
  wire [255:0] _data_io_dinb_T_2 = {dp_write_line_3,dp_write_line_2,dp_write_line_1,dp_write_line_0}; // @[Dcache.scala 187:113]
  wire  _meta_io_update_T_2 = wb_valid ? 1'h0 : _data_io_web_T_1; // @[Dcache.scala 195:30]
  wire [63:0] _io_bar_req_data_T = dp_mmio_valid ? dp_mmio_req_wdata : io_cpu_req_bits_wdata; // @[Dcache.scala 205:55]
  wire [31:0] _io_bar_req_addr_T_1 = _T_22 ? wb_dirty_addr : wb_refill_addr; // @[Dcache.scala 206:40]
  wire [31:0] _io_bar_req_addr_T_2 = dp_mmio_valid ? dp_mmio_req_addr : io_cpu_req_bits_addr; // @[Dcache.scala 206:106]
  wire [2:0] _io_bar_req_mtype_T = dp_mmio_valid ? dp_mmio_req_mtype : io_cpu_req_bits_mtype; // @[Dcache.scala 207:52]
  wire  _io_bar_req_valid_T_3 = dp_mmio_valid ? _dp_mmio_stall_T : df_mmio_valid; // @[Dcache.scala 209:72]
  wire  _io_bar_req_wen_T_1 = dp_mmio_valid ? dp_mmio_req_wen : io_cpu_req_bits_wen; // @[Dcache.scala 213:70]
  wire  _wb_state_T = meta_io_dirty ? 1'h0 : 1'h1; // @[Dcache.scala 220:26]
  wire [31:0] _wb_dirty_addr_T = {meta_io_tag_fetch,dp_index,5'h0}; // @[Cat.scala 30:58]
  wire [255:0] _wb_dirty_data_T = {dp_fetch_line_3,dp_fetch_line_2,dp_fetch_line_1,dp_fetch_line_0}; // @[Dcache.scala 222:43]
  wire  _GEN_28 = _dp_index_T ? _wb_state_T : wb_state; // @[Dcache.scala 219:20 Dcache.scala 220:20 Dcache.scala 201:25]
  wire  _GEN_52 = wb_state | _meta_io_update_T_2; // @[Conditional.scala 39:67 Dcache.scala 243:24 Dcache.scala 195:24]
  wire  _GEN_55 = _T_22 ? _meta_io_update_T_2 : _GEN_52; // @[Conditional.scala 40:58 Dcache.scala 195:24]
  DualPortBRAM_2 data ( // @[Dcache.scala 66:20]
    .clock(data_clock),
    .reset(data_reset),
    .io_web(data_io_web),
    .io_addra(data_io_addra),
    .io_addrb(data_io_addrb),
    .io_dinb(data_io_dinb),
    .io_douta(data_io_douta)
  );
  MetaDataBRAM meta ( // @[Dcache.scala 67:20]
    .clock(meta_clock),
    .reset(meta_reset),
    .io_index_fetch(meta_io_index_fetch),
    .io_index_update(meta_io_index_update),
    .io_tag_update(meta_io_tag_update),
    .io_update(meta_io_update),
    .io_write(meta_io_write),
    .io_hit(meta_io_hit),
    .io_tag_fetch(meta_io_tag_fetch),
    .io_dirty(meta_io_dirty)
  );
  assign io_cpu_resp_valid = wb_resp_valid | dp_resp_valid | dp_mmio_resp_valid; // @[Dcache.scala 179:63]
  assign io_cpu_resp_bits_rdata_0 = _T_13[31:0]; // @[Dcache.scala 184:42]
  assign io_cpu_resp_bits_rdata_1 = _T_13[63:32]; // @[Dcache.scala 184:42]
  assign io_bar_req_valid = wb_valid ? wb_valid & _dp_mmio_stall_T : _io_bar_req_valid_T_3; // @[Dcache.scala 209:26]
  assign io_bar_req_wen = wb_valid ? _T_22 : _io_bar_req_wen_T_1; // @[Dcache.scala 213:26]
  assign io_bar_req_addr = wb_valid ? _io_bar_req_addr_T_1 : _io_bar_req_addr_T_2; // @[Dcache.scala 206:26]
  assign io_bar_req_data = wb_valid ? wb_dirty_data : {{192'd0}, _io_bar_req_data_T}; // @[Dcache.scala 205:26]
  assign io_bar_req_mtype = wb_valid ? 3'h4 : _io_bar_req_mtype_T; // @[Dcache.scala 207:26]
  assign data_clock = clock;
  assign data_reset = reset;
  assign data_io_web = wb_valid ? wb_write_cache : dp_resp_valid & dp_req_wen; // @[Dcache.scala 186:23]
  assign data_io_addra = io_cpu_req_bits_addr[13:5]; // @[Dcache.scala 74:49]
  assign data_io_addrb = wb_valid ? wb_index : dp_index; // @[Dcache.scala 189:23]
  assign data_io_dinb = wb_valid ? _data_io_dinb_T_1 : _data_io_dinb_T_2; // @[Dcache.scala 187:23]
  assign meta_clock = clock;
  assign meta_reset = reset;
  assign meta_io_index_fetch = io_cpu_req_bits_addr[13:5]; // @[Dcache.scala 74:49]
  assign meta_io_index_update = wb_valid ? wb_index : dp_index; // @[Dcache.scala 193:30]
  assign meta_io_tag_update = wb_valid ? wb_tag : dp_tag; // @[Dcache.scala 192:30]
  assign meta_io_update = wb_valid ? _GEN_55 : _meta_io_update_T_2; // @[Dcache.scala 237:19 Dcache.scala 195:24]
  assign meta_io_write = wb_valid ? wb_req_wen : dp_req_wen; // @[Dcache.scala 194:30]
  always @(posedge clock) begin
    if (reset) begin // @[Dcache.scala 97:31]
      wb_valid <= 1'h0; // @[Dcache.scala 97:31]
    end else if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_valid <= _dp_valid_T_1; // @[Dcache.scala 223:20]
    end
    if (reset) begin // @[Dcache.scala 201:25]
      wb_state <= 1'h0; // @[Dcache.scala 201:25]
    end else if (wb_valid) begin // @[Dcache.scala 237:19]
      if (_T_22) begin // @[Conditional.scala 40:58]
        wb_state <= io_bar_resp_valid | wb_state; // @[Dcache.scala 240:18]
      end else begin
        wb_state <= _GEN_28;
      end
    end else begin
      wb_state <= _GEN_28;
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_index <= df_index; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_tag <= df_tag; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_offset <= df_offset; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_req_addr <= io_cpu_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_req_wdata <= io_cpu_req_bits_wdata; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_req_wen <= io_cpu_req_bits_wen; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Reg.scala 16:19]
      dp_req_mtype <= io_cpu_req_bits_mtype; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Dcache.scala 87:36]
      dp_valid <= 1'h0; // @[Dcache.scala 87:36]
    end else if (dp_valid & ~meta_io_hit | wb_stall | df_mmio_valid | dp_mmio_stall) begin // @[Dcache.scala 157:23]
      dp_valid <= 1'h0;
    end else begin
      dp_valid <= io_cpu_req_valid;
    end
    if (_dp_mmio_valid_T) begin // @[Reg.scala 16:19]
      dp_mmio_valid <= df_mmio_valid; // @[Reg.scala 16:23]
    end
    if (_dp_mmio_valid_T) begin // @[Reg.scala 16:19]
      dp_mmio_req_addr <= io_cpu_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_dp_mmio_valid_T) begin // @[Reg.scala 16:19]
      dp_mmio_req_wdata <= io_cpu_req_bits_wdata; // @[Reg.scala 16:23]
    end
    if (_dp_mmio_valid_T) begin // @[Reg.scala 16:19]
      dp_mmio_req_wen <= io_cpu_req_bits_wen; // @[Reg.scala 16:23]
    end
    if (_dp_mmio_valid_T) begin // @[Reg.scala 16:19]
      dp_mmio_req_mtype <= io_cpu_req_bits_mtype; // @[Reg.scala 16:23]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_dirty_data <= _wb_dirty_data_T; // @[Dcache.scala 222:20]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_dirty_addr <= _wb_dirty_addr_T; // @[Dcache.scala 221:20]
    end
    if (reset) begin // @[Dcache.scala 99:31]
      wb_req_wdata <= 64'h0; // @[Dcache.scala 99:31]
    end else if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_req_wdata <= dp_req_wdata; // @[Dcache.scala 225:20]
    end
    if (reset) begin // @[Dcache.scala 99:31]
      wb_req_wen <= 1'h0; // @[Dcache.scala 99:31]
    end else if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_req_wen <= dp_req_wen; // @[Dcache.scala 225:20]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_index <= dp_index; // @[Dcache.scala 226:20]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_tag <= dp_tag; // @[Dcache.scala 227:20]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_offset <= {{3'd0}, dp_offset}; // @[Dcache.scala 228:20]
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      if (3'h2 == dp_req_mtype) begin // @[Mux.scala 80:57]
        wb_mask <= 64'hffffffff;
      end else if (3'h0 == dp_req_mtype) begin // @[Mux.scala 80:57]
        wb_mask <= 64'hff;
      end else if (3'h1 == dp_req_mtype) begin // @[Mux.scala 80:57]
        wb_mask <= 64'hffff;
      end else begin
        wb_mask <= 64'hffffffffffffffff;
      end
    end
    if (_dp_index_T) begin // @[Dcache.scala 219:20]
      wb_shift <= dp_shift; // @[Dcache.scala 230:20]
    end
    REG <= data_io_web & data_io_addra == data_io_addrb; // @[Dcache.scala 153:44]
    REG_1_0 <= _WIRE_1[63:0]; // @[Dcache.scala 154:34]
    REG_1_1 <= _WIRE_1[127:64]; // @[Dcache.scala 154:34]
    REG_1_2 <= _WIRE_1[191:128]; // @[Dcache.scala 154:34]
    REG_1_3 <= _WIRE_1[255:192]; // @[Dcache.scala 154:34]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_state = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dp_index = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  dp_tag = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  dp_offset = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  dp_req_addr = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  dp_req_wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  dp_req_wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dp_req_mtype = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  dp_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dp_mmio_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dp_mmio_req_addr = _RAND_11[31:0];
  _RAND_12 = {2{`RANDOM}};
  dp_mmio_req_wdata = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  dp_mmio_req_wen = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dp_mmio_req_mtype = _RAND_14[2:0];
  _RAND_15 = {8{`RANDOM}};
  wb_dirty_data = _RAND_15[255:0];
  _RAND_16 = {1{`RANDOM}};
  wb_dirty_addr = _RAND_16[31:0];
  _RAND_17 = {2{`RANDOM}};
  wb_req_wdata = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  wb_req_wen = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  wb_index = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  wb_tag = _RAND_20[17:0];
  _RAND_21 = {1{`RANDOM}};
  wb_offset = _RAND_21[4:0];
  _RAND_22 = {2{`RANDOM}};
  wb_mask = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  wb_shift = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  REG = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  REG_1_0 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  REG_1_1 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  REG_1_2 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  REG_1_3 = _RAND_28[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DcacheDPFilter(
  input          clock,
  input          reset,
  input          io_dcache_cpu_req_valid,
  input  [31:0]  io_dcache_cpu_req_bits_addr,
  input  [63:0]  io_dcache_cpu_req_bits_wdata,
  input          io_dcache_cpu_req_bits_wen,
  input  [2:0]   io_dcache_cpu_req_bits_mtype,
  output         io_dcache_cpu_resp_valid,
  output [31:0]  io_dcache_cpu_resp_bits_rdata_0,
  output [31:0]  io_dcache_cpu_resp_bits_rdata_1,
  output         io_dcache_bar_req_valid,
  output         io_dcache_bar_req_wen,
  output [31:0]  io_dcache_bar_req_addr,
  output [255:0] io_dcache_bar_req_data,
  output [2:0]   io_dcache_bar_req_mtype,
  input          io_dcache_bar_resp_valid,
  input  [255:0] io_dcache_bar_resp_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  dcache_clock; // @[Dcache.scala 260:22]
  wire  dcache_reset; // @[Dcache.scala 260:22]
  wire  dcache_io_cpu_req_valid; // @[Dcache.scala 260:22]
  wire [31:0] dcache_io_cpu_req_bits_addr; // @[Dcache.scala 260:22]
  wire [63:0] dcache_io_cpu_req_bits_wdata; // @[Dcache.scala 260:22]
  wire  dcache_io_cpu_req_bits_wen; // @[Dcache.scala 260:22]
  wire [2:0] dcache_io_cpu_req_bits_mtype; // @[Dcache.scala 260:22]
  wire  dcache_io_cpu_resp_valid; // @[Dcache.scala 260:22]
  wire [31:0] dcache_io_cpu_resp_bits_rdata_0; // @[Dcache.scala 260:22]
  wire [31:0] dcache_io_cpu_resp_bits_rdata_1; // @[Dcache.scala 260:22]
  wire  dcache_io_bar_req_valid; // @[Dcache.scala 260:22]
  wire  dcache_io_bar_req_wen; // @[Dcache.scala 260:22]
  wire [31:0] dcache_io_bar_req_addr; // @[Dcache.scala 260:22]
  wire [255:0] dcache_io_bar_req_data; // @[Dcache.scala 260:22]
  wire [2:0] dcache_io_bar_req_mtype; // @[Dcache.scala 260:22]
  wire  dcache_io_bar_resp_valid; // @[Dcache.scala 260:22]
  wire [255:0] dcache_io_bar_resp_data; // @[Dcache.scala 260:22]
  reg [63:0] mtime; // @[Dcache.scala 265:20]
  reg [63:0] mtimecmp; // @[Dcache.scala 266:23]
  reg  counter; // @[Dcache.scala 267:26]
  wire [5:0] _GEN_15 = {{5'd0}, counter}; // @[Dcache.scala 269:28]
  wire  _counter_T = _GEN_15 == 6'h32; // @[Dcache.scala 269:28]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[Dcache.scala 271:22]
  wire [63:0] _GEN_0 = _counter_T ? _mtime_T_1 : mtime; // @[Dcache.scala 270:36 Dcache.scala 271:13 Dcache.scala 265:20]
  wire  _hit_clint_addr_T = io_dcache_cpu_req_bits_addr == 32'h200bff8; // @[Dcache.scala 280:54]
  wire  _hit_clint_addr_T_1 = io_dcache_cpu_req_bits_addr == 32'h2004000; // @[Dcache.scala 280:102]
  wire  hit_clint_addr = io_dcache_cpu_req_bits_addr == 32'h200bff8 | io_dcache_cpu_req_bits_addr == 32'h2004000; // @[Dcache.scala 280:71]
  reg [31:0] last_req_addr; // @[Dcache.scala 281:33]
  reg  io_dcache_cpu_resp_valid_REG; // @[Dcache.scala 298:42]
  reg  io_dcache_cpu_resp_valid_REG_1; // @[Dcache.scala 302:42]
  wire [31:0] _GEN_9 = last_req_addr == 32'h2004000 ? mtimecmp[31:0] : dcache_io_cpu_resp_bits_rdata_0; // @[Dcache.scala 299:52 Dcache.scala 300:40 Dcache.scala 262:13]
  wire [31:0] _GEN_10 = last_req_addr == 32'h2004000 ? mtimecmp[63:32] : dcache_io_cpu_resp_bits_rdata_1; // @[Dcache.scala 299:52 Dcache.scala 301:40 Dcache.scala 262:13]
  wire  _GEN_11 = last_req_addr == 32'h2004000 ? io_dcache_cpu_resp_valid_REG_1 : dcache_io_cpu_resp_valid; // @[Dcache.scala 299:52 Dcache.scala 302:32 Dcache.scala 262:13]
  DcacheDP dcache ( // @[Dcache.scala 260:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_wdata(dcache_io_cpu_req_bits_wdata),
    .io_cpu_req_bits_wen(dcache_io_cpu_req_bits_wen),
    .io_cpu_req_bits_mtype(dcache_io_cpu_req_bits_mtype),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_rdata_0(dcache_io_cpu_resp_bits_rdata_0),
    .io_cpu_resp_bits_rdata_1(dcache_io_cpu_resp_bits_rdata_1),
    .io_bar_req_valid(dcache_io_bar_req_valid),
    .io_bar_req_wen(dcache_io_bar_req_wen),
    .io_bar_req_addr(dcache_io_bar_req_addr),
    .io_bar_req_data(dcache_io_bar_req_data),
    .io_bar_req_mtype(dcache_io_bar_req_mtype),
    .io_bar_resp_valid(dcache_io_bar_resp_valid),
    .io_bar_resp_data(dcache_io_bar_resp_data)
  );
  assign io_dcache_cpu_resp_valid = last_req_addr == 32'h200bff8 ? io_dcache_cpu_resp_valid_REG : _GEN_11; // @[Dcache.scala 295:43 Dcache.scala 298:32]
  assign io_dcache_cpu_resp_bits_rdata_0 = last_req_addr == 32'h200bff8 ? mtime[31:0] : _GEN_9; // @[Dcache.scala 295:43 Dcache.scala 296:40]
  assign io_dcache_cpu_resp_bits_rdata_1 = last_req_addr == 32'h200bff8 ? mtime[63:32] : _GEN_10; // @[Dcache.scala 295:43 Dcache.scala 297:40]
  assign io_dcache_bar_req_valid = dcache_io_bar_req_valid; // @[Dcache.scala 262:13]
  assign io_dcache_bar_req_wen = dcache_io_bar_req_wen; // @[Dcache.scala 262:13]
  assign io_dcache_bar_req_addr = dcache_io_bar_req_addr; // @[Dcache.scala 262:13]
  assign io_dcache_bar_req_data = dcache_io_bar_req_data; // @[Dcache.scala 262:13]
  assign io_dcache_bar_req_mtype = dcache_io_bar_req_mtype; // @[Dcache.scala 262:13]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_req_valid = hit_clint_addr ? 1'h0 : io_dcache_cpu_req_valid; // @[Dcache.scala 282:27 Dcache.scala 283:31 Dcache.scala 262:13]
  assign dcache_io_cpu_req_bits_addr = io_dcache_cpu_req_bits_addr; // @[Dcache.scala 262:13]
  assign dcache_io_cpu_req_bits_wdata = io_dcache_cpu_req_bits_wdata; // @[Dcache.scala 262:13]
  assign dcache_io_cpu_req_bits_wen = io_dcache_cpu_req_bits_wen; // @[Dcache.scala 262:13]
  assign dcache_io_cpu_req_bits_mtype = io_dcache_cpu_req_bits_mtype; // @[Dcache.scala 262:13]
  assign dcache_io_bar_resp_valid = io_dcache_bar_resp_valid; // @[Dcache.scala 262:13]
  assign dcache_io_bar_resp_data = io_dcache_bar_resp_data; // @[Dcache.scala 262:13]
  always @(posedge clock) begin
    if (hit_clint_addr) begin // @[Dcache.scala 282:27]
      if (io_dcache_cpu_req_valid & io_dcache_cpu_req_bits_wen) begin // @[Dcache.scala 285:68]
        if (_hit_clint_addr_T) begin // @[Dcache.scala 286:61]
          mtime <= io_dcache_cpu_req_bits_wdata; // @[Dcache.scala 287:17]
        end else begin
          mtime <= _GEN_0;
        end
      end else begin
        mtime <= _GEN_0;
      end
    end else begin
      mtime <= _GEN_0;
    end
    if (hit_clint_addr) begin // @[Dcache.scala 282:27]
      if (io_dcache_cpu_req_valid & io_dcache_cpu_req_bits_wen) begin // @[Dcache.scala 285:68]
        if (!(_hit_clint_addr_T)) begin // @[Dcache.scala 286:61]
          if (_hit_clint_addr_T_1) begin // @[Dcache.scala 288:70]
            mtimecmp <= io_dcache_cpu_req_bits_wdata; // @[Dcache.scala 289:20]
          end
        end
      end
    end
    if (reset) begin // @[Dcache.scala 267:26]
      counter <= 1'h0; // @[Dcache.scala 267:26]
    end else if (_GEN_15 == 6'h32) begin // @[Dcache.scala 269:19]
      counter <= 1'h0;
    end else begin
      counter <= counter + 1'h1;
    end
    last_req_addr <= io_dcache_cpu_req_bits_addr; // @[Dcache.scala 281:33]
    io_dcache_cpu_resp_valid_REG <= io_dcache_cpu_req_valid; // @[Dcache.scala 298:42]
    io_dcache_cpu_resp_valid_REG_1 <= io_dcache_cpu_req_valid; // @[Dcache.scala 302:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  last_req_addr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  io_dcache_cpu_resp_valid_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_dcache_cpu_resp_valid_REG_1 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimMem(
  input          clock,
  input          reset,
  input          io_icache_io_req_valid,
  input  [31:0]  io_icache_io_req_addr,
  output         io_icache_io_resp_valid,
  output [255:0] io_icache_io_resp_data,
  input          io_dcache_io_req_valid,
  input          io_dcache_io_req_wen,
  input  [31:0]  io_dcache_io_req_addr,
  input  [255:0] io_dcache_io_req_data,
  input  [2:0]   io_dcache_io_req_mtype,
  output         io_dcache_io_resp_valid,
  output [255:0] io_dcache_io_resp_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [255:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] memory [0:67108863]; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_0_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_0_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_0_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_0_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_1_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_1_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_1_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_1_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_2_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_2_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_2_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_2_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_3_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_3_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_3_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_3_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_4_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_4_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_4_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_4_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_5_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_5_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_5_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_5_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_6_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_6_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_6_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_6_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_7_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_7_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_7_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_7_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_8_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_8_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_8_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_8_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_9_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_9_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_9_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_9_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_10_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_10_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_10_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_10_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_11_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_11_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_11_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_11_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_12_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_12_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_12_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_12_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_13_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_13_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_13_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_13_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_14_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_14_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_14_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_14_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_15_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_15_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_15_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_15_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_16_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_16_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_16_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_16_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_17_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_17_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_17_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_17_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_18_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_18_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_18_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_18_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_19_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_19_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_19_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_19_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_20_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_20_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_20_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_20_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_21_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_21_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_21_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_21_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_22_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_22_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_22_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_22_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_23_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_23_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_23_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_23_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_24_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_24_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_24_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_24_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_25_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_25_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_25_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_25_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_26_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_26_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_26_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_26_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_27_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_27_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_27_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_27_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_28_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_28_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_28_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_28_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_29_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_29_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_29_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_29_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_30_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_30_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_30_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_30_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_icandidates_31_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_icandidates_31_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_dcandidates_31_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_dcandidates_31_MPORT_addr; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_1_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_1_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_1_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_1_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_2_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_2_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_2_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_2_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_3_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_3_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_3_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_3_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_4_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_4_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_4_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_4_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_5_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_5_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_5_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_5_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_6_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_6_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_6_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_6_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_7_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_7_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_7_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_7_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_8_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_8_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_8_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_8_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_9_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_9_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_9_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_9_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_10_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_10_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_10_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_10_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_11_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_11_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_11_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_11_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_12_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_12_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_12_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_12_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_13_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_13_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_13_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_13_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_14_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_14_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_14_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_14_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_15_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_15_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_15_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_15_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_16_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_16_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_16_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_16_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_17_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_17_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_17_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_17_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_18_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_18_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_18_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_18_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_19_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_19_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_19_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_19_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_20_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_20_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_20_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_20_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_21_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_21_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_21_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_21_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_22_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_22_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_22_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_22_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_23_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_23_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_23_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_23_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_24_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_24_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_24_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_24_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_25_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_25_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_25_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_25_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_26_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_26_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_26_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_26_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_27_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_27_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_27_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_27_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_28_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_28_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_28_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_28_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_29_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_29_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_29_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_29_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_30_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_30_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_30_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_30_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_31_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_31_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_31_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_31_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_32_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_32_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_32_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_32_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_33_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_33_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_33_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_33_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_34_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_34_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_34_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_34_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_35_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_35_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_35_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_35_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_36_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_36_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_36_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_36_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_37_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_37_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_37_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_37_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_38_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_38_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_38_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_38_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_39_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_39_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_39_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_39_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_40_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_40_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_40_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_40_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_41_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_41_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_41_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_41_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_42_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_42_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_42_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_42_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_43_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_43_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_43_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_43_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_44_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_44_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_44_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_44_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_45_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_45_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_45_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_45_en; // @[SimMem.scala 42:19]
  wire [7:0] memory_MPORT_46_data; // @[SimMem.scala 42:19]
  wire [25:0] memory_MPORT_46_addr; // @[SimMem.scala 42:19]
  wire  memory_MPORT_46_mask; // @[SimMem.scala 42:19]
  wire  memory_MPORT_46_en; // @[SimMem.scala 42:19]
  wire  _GEN_0 = io_dcache_io_req_addr[29:0] >= 30'h4000000 ? 1'h0 : 1'h1; // @[SimMem.scala 25:56 SimMem.scala 26:17]
  wire  _T_6 = io_dcache_io_req_addr == 32'h10000000 & io_dcache_io_req_wen & ~io_dcache_io_resp_valid; // @[SimMem.scala 29:83]
  wire  _T_9 = ~reset; // @[SimMem.scala 30:14]
  wire  write_ram = io_dcache_io_req_valid ? _GEN_0 : 1'h1; // @[SimMem.scala 24:32]
  wire  _T_10 = io_icache_io_req_addr >= 32'h84000000; // @[SimMem.scala 35:32]
  wire [32:0] _icandidates_0_T = {{1'd0}, io_icache_io_req_addr}; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_0_T_2 = 32'h3ffffff & _icandidates_0_T[31:0]; // @[SimMem.scala 46:44]
  wire [29:0] dcandidates_0_hi = io_dcache_io_req_addr[31:2]; // @[SimMem.scala 47:72]
  wire [31:0] _dcandidates_0_T = {dcandidates_0_hi,2'h0}; // @[Cat.scala 30:58]
  wire [32:0] _dcandidates_0_T_1 = {{1'd0}, _dcandidates_0_T}; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_0_T_3 = 32'h3ffffff & _dcandidates_0_T_1[31:0]; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_1_T_1 = io_icache_io_req_addr + 32'h1; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_1_T_2 = 32'h3ffffff & _icandidates_1_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_1_T_2 = _dcandidates_0_T + 32'h1; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_1_T_3 = 32'h3ffffff & _dcandidates_1_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_2_T_1 = io_icache_io_req_addr + 32'h2; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_2_T_2 = 32'h3ffffff & _icandidates_2_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_2_T_2 = _dcandidates_0_T + 32'h2; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_2_T_3 = 32'h3ffffff & _dcandidates_2_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_3_T_1 = io_icache_io_req_addr + 32'h3; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_3_T_2 = 32'h3ffffff & _icandidates_3_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_3_T_2 = _dcandidates_0_T + 32'h3; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_3_T_3 = 32'h3ffffff & _dcandidates_3_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_4_T_1 = io_icache_io_req_addr + 32'h4; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_4_T_2 = 32'h3ffffff & _icandidates_4_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_4_T_2 = _dcandidates_0_T + 32'h4; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_4_T_3 = 32'h3ffffff & _dcandidates_4_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_5_T_1 = io_icache_io_req_addr + 32'h5; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_5_T_2 = 32'h3ffffff & _icandidates_5_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_5_T_2 = _dcandidates_0_T + 32'h5; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_5_T_3 = 32'h3ffffff & _dcandidates_5_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_6_T_1 = io_icache_io_req_addr + 32'h6; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_6_T_2 = 32'h3ffffff & _icandidates_6_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_6_T_2 = _dcandidates_0_T + 32'h6; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_6_T_3 = 32'h3ffffff & _dcandidates_6_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_7_T_1 = io_icache_io_req_addr + 32'h7; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_7_T_2 = 32'h3ffffff & _icandidates_7_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_7_T_2 = _dcandidates_0_T + 32'h7; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_7_T_3 = 32'h3ffffff & _dcandidates_7_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_8_T_1 = io_icache_io_req_addr + 32'h8; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_8_T_2 = 32'h3ffffff & _icandidates_8_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_8_T_2 = _dcandidates_0_T + 32'h8; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_8_T_3 = 32'h3ffffff & _dcandidates_8_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_9_T_1 = io_icache_io_req_addr + 32'h9; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_9_T_2 = 32'h3ffffff & _icandidates_9_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_9_T_2 = _dcandidates_0_T + 32'h9; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_9_T_3 = 32'h3ffffff & _dcandidates_9_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_10_T_1 = io_icache_io_req_addr + 32'ha; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_10_T_2 = 32'h3ffffff & _icandidates_10_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_10_T_2 = _dcandidates_0_T + 32'ha; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_10_T_3 = 32'h3ffffff & _dcandidates_10_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_11_T_1 = io_icache_io_req_addr + 32'hb; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_11_T_2 = 32'h3ffffff & _icandidates_11_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_11_T_2 = _dcandidates_0_T + 32'hb; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_11_T_3 = 32'h3ffffff & _dcandidates_11_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_12_T_1 = io_icache_io_req_addr + 32'hc; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_12_T_2 = 32'h3ffffff & _icandidates_12_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_12_T_2 = _dcandidates_0_T + 32'hc; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_12_T_3 = 32'h3ffffff & _dcandidates_12_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_13_T_1 = io_icache_io_req_addr + 32'hd; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_13_T_2 = 32'h3ffffff & _icandidates_13_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_13_T_2 = _dcandidates_0_T + 32'hd; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_13_T_3 = 32'h3ffffff & _dcandidates_13_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_14_T_1 = io_icache_io_req_addr + 32'he; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_14_T_2 = 32'h3ffffff & _icandidates_14_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_14_T_2 = _dcandidates_0_T + 32'he; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_14_T_3 = 32'h3ffffff & _dcandidates_14_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_15_T_1 = io_icache_io_req_addr + 32'hf; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_15_T_2 = 32'h3ffffff & _icandidates_15_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_15_T_2 = _dcandidates_0_T + 32'hf; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_15_T_3 = 32'h3ffffff & _dcandidates_15_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_16_T_1 = io_icache_io_req_addr + 32'h10; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_16_T_2 = 32'h3ffffff & _icandidates_16_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_16_T_2 = _dcandidates_0_T + 32'h10; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_16_T_3 = 32'h3ffffff & _dcandidates_16_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_17_T_1 = io_icache_io_req_addr + 32'h11; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_17_T_2 = 32'h3ffffff & _icandidates_17_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_17_T_2 = _dcandidates_0_T + 32'h11; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_17_T_3 = 32'h3ffffff & _dcandidates_17_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_18_T_1 = io_icache_io_req_addr + 32'h12; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_18_T_2 = 32'h3ffffff & _icandidates_18_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_18_T_2 = _dcandidates_0_T + 32'h12; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_18_T_3 = 32'h3ffffff & _dcandidates_18_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_19_T_1 = io_icache_io_req_addr + 32'h13; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_19_T_2 = 32'h3ffffff & _icandidates_19_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_19_T_2 = _dcandidates_0_T + 32'h13; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_19_T_3 = 32'h3ffffff & _dcandidates_19_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_20_T_1 = io_icache_io_req_addr + 32'h14; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_20_T_2 = 32'h3ffffff & _icandidates_20_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_20_T_2 = _dcandidates_0_T + 32'h14; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_20_T_3 = 32'h3ffffff & _dcandidates_20_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_21_T_1 = io_icache_io_req_addr + 32'h15; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_21_T_2 = 32'h3ffffff & _icandidates_21_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_21_T_2 = _dcandidates_0_T + 32'h15; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_21_T_3 = 32'h3ffffff & _dcandidates_21_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_22_T_1 = io_icache_io_req_addr + 32'h16; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_22_T_2 = 32'h3ffffff & _icandidates_22_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_22_T_2 = _dcandidates_0_T + 32'h16; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_22_T_3 = 32'h3ffffff & _dcandidates_22_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_23_T_1 = io_icache_io_req_addr + 32'h17; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_23_T_2 = 32'h3ffffff & _icandidates_23_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_23_T_2 = _dcandidates_0_T + 32'h17; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_23_T_3 = 32'h3ffffff & _dcandidates_23_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_24_T_1 = io_icache_io_req_addr + 32'h18; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_24_T_2 = 32'h3ffffff & _icandidates_24_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_24_T_2 = _dcandidates_0_T + 32'h18; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_24_T_3 = 32'h3ffffff & _dcandidates_24_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_25_T_1 = io_icache_io_req_addr + 32'h19; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_25_T_2 = 32'h3ffffff & _icandidates_25_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_25_T_2 = _dcandidates_0_T + 32'h19; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_25_T_3 = 32'h3ffffff & _dcandidates_25_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_26_T_1 = io_icache_io_req_addr + 32'h1a; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_26_T_2 = 32'h3ffffff & _icandidates_26_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_26_T_2 = _dcandidates_0_T + 32'h1a; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_26_T_3 = 32'h3ffffff & _dcandidates_26_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_27_T_1 = io_icache_io_req_addr + 32'h1b; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_27_T_2 = 32'h3ffffff & _icandidates_27_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_27_T_2 = _dcandidates_0_T + 32'h1b; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_27_T_3 = 32'h3ffffff & _dcandidates_27_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_28_T_1 = io_icache_io_req_addr + 32'h1c; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_28_T_2 = 32'h3ffffff & _icandidates_28_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_28_T_2 = _dcandidates_0_T + 32'h1c; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_28_T_3 = 32'h3ffffff & _dcandidates_28_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_29_T_1 = io_icache_io_req_addr + 32'h1d; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_29_T_2 = 32'h3ffffff & _icandidates_29_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_29_T_2 = _dcandidates_0_T + 32'h1d; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_29_T_3 = 32'h3ffffff & _dcandidates_29_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_30_T_1 = io_icache_io_req_addr + 32'h1e; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_30_T_2 = 32'h3ffffff & _icandidates_30_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_30_T_2 = _dcandidates_0_T + 32'h1e; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_30_T_3 = 32'h3ffffff & _dcandidates_30_T_2; // @[SimMem.scala 47:44]
  wire [31:0] _icandidates_31_T_1 = io_icache_io_req_addr + 32'h1f; // @[SimMem.scala 46:69]
  wire [31:0] _icandidates_31_T_2 = 32'h3ffffff & _icandidates_31_T_1; // @[SimMem.scala 46:44]
  wire [31:0] _dcandidates_31_T_2 = _dcandidates_0_T + 32'h1f; // @[SimMem.scala 47:89]
  wire [31:0] _dcandidates_31_T_3 = 32'h3ffffff & _dcandidates_31_T_2; // @[SimMem.scala 47:44]
  wire [7:0] dcandidates_0 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_0_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_1 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_1_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_2 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_2_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_3 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_3_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_4 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_4_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_5 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_5_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_6 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_6_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_7 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_7_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_8 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_8_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_9 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_9_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_10 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_10_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_11 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_11_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_12 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_12_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_13 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_13_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_14 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_14_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_15 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_15_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_16 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_16_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_17 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_17_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_18 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_18_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_19 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_19_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_20 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_20_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_21 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_21_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_22 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_22_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_23 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_23_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_24 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_24_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_25 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_25_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_26 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_26_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_27 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_27_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_28 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_28_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_29 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_29_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_30 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_30_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  wire [7:0] dcandidates_31 = io_dcache_io_req_valid & io_dcache_io_req_addr == 32'h10000003 ? 8'h0 :
    memory_dcandidates_31_MPORT_data; // @[SimMem.scala 57:78 SimMem.scala 58:17 SimMem.scala 47:20]
  reg  io_icache_io_resp_valid_REG; // @[SimMem.scala 63:37]
  wire [7:0] icandidates_1 = memory_icandidates_1_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_0 = memory_icandidates_0_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_3 = memory_icandidates_3_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_2 = memory_icandidates_2_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_5 = memory_icandidates_5_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_4 = memory_icandidates_4_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_7 = memory_icandidates_7_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_6 = memory_icandidates_6_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [63:0] io_icache_io_resp_data_lo_lo = {icandidates_7,icandidates_6,icandidates_5,icandidates_4,icandidates_3,
    icandidates_2,icandidates_1,icandidates_0}; // @[SimMem.scala 64:50]
  wire [7:0] icandidates_9 = memory_icandidates_9_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_8 = memory_icandidates_8_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_11 = memory_icandidates_11_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_10 = memory_icandidates_10_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_13 = memory_icandidates_13_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_12 = memory_icandidates_12_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_15 = memory_icandidates_15_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_14 = memory_icandidates_14_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [127:0] io_icache_io_resp_data_lo = {icandidates_15,icandidates_14,icandidates_13,icandidates_12,icandidates_11,
    icandidates_10,icandidates_9,icandidates_8,io_icache_io_resp_data_lo_lo}; // @[SimMem.scala 64:50]
  wire [7:0] icandidates_17 = memory_icandidates_17_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_16 = memory_icandidates_16_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_19 = memory_icandidates_19_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_18 = memory_icandidates_18_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_21 = memory_icandidates_21_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_20 = memory_icandidates_20_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_23 = memory_icandidates_23_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_22 = memory_icandidates_22_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [63:0] io_icache_io_resp_data_hi_lo = {icandidates_23,icandidates_22,icandidates_21,icandidates_20,icandidates_19
    ,icandidates_18,icandidates_17,icandidates_16}; // @[SimMem.scala 64:50]
  wire [7:0] icandidates_25 = memory_icandidates_25_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_24 = memory_icandidates_24_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_27 = memory_icandidates_27_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_26 = memory_icandidates_26_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_29 = memory_icandidates_29_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_28 = memory_icandidates_28_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_31 = memory_icandidates_31_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [7:0] icandidates_30 = memory_icandidates_30_MPORT_data; // @[SimMem.scala 20:25 SimMem.scala 46:20]
  wire [127:0] io_icache_io_resp_data_hi = {icandidates_31,icandidates_30,icandidates_29,icandidates_28,icandidates_27,
    icandidates_26,icandidates_25,icandidates_24,io_icache_io_resp_data_hi_lo}; // @[SimMem.scala 64:50]
  reg [255:0] io_icache_io_resp_data_REG; // @[SimMem.scala 64:37]
  reg  io_dcache_io_resp_valid_REG; // @[SimMem.scala 65:37]
  wire [63:0] io_dcache_io_resp_data_lo_lo = {dcandidates_7,dcandidates_6,dcandidates_5,dcandidates_4,dcandidates_3,
    dcandidates_2,dcandidates_1,dcandidates_0}; // @[SimMem.scala 66:50]
  wire [127:0] io_dcache_io_resp_data_lo = {dcandidates_15,dcandidates_14,dcandidates_13,dcandidates_12,dcandidates_11,
    dcandidates_10,dcandidates_9,dcandidates_8,io_dcache_io_resp_data_lo_lo}; // @[SimMem.scala 66:50]
  wire [63:0] io_dcache_io_resp_data_hi_lo = {dcandidates_23,dcandidates_22,dcandidates_21,dcandidates_20,dcandidates_19
    ,dcandidates_18,dcandidates_17,dcandidates_16}; // @[SimMem.scala 66:50]
  wire [127:0] io_dcache_io_resp_data_hi = {dcandidates_31,dcandidates_30,dcandidates_29,dcandidates_28,dcandidates_27,
    dcandidates_26,dcandidates_25,dcandidates_24,io_dcache_io_resp_data_hi_lo}; // @[SimMem.scala 66:50]
  reg [255:0] io_dcache_io_resp_data_REG; // @[SimMem.scala 66:37]
  wire  _T_16 = io_dcache_io_req_wen & write_ram & io_dcache_io_req_valid; // @[SimMem.scala 70:42]
  wire  _T_17 = 3'h0 == io_dcache_io_req_mtype; // @[Conditional.scala 37:30]
  wire [31:0] _T_18 = io_dcache_io_req_addr & 32'h3ffffff; // @[SimMem.scala 74:44]
  wire  _T_21 = 3'h1 == io_dcache_io_req_mtype; // @[Conditional.scala 37:30]
  wire [31:0] _T_26 = io_dcache_io_req_addr + 32'h1; // @[SimMem.scala 79:45]
  wire [31:0] _T_27 = _T_26 & 32'h3ffffff; // @[SimMem.scala 79:52]
  wire  _T_30 = 3'h2 == io_dcache_io_req_mtype; // @[Conditional.scala 37:30]
  wire [31:0] _T_40 = io_dcache_io_req_addr + 32'h2; // @[SimMem.scala 85:45]
  wire [31:0] _T_41 = _T_40 & 32'h3ffffff; // @[SimMem.scala 85:52]
  wire [31:0] _T_45 = io_dcache_io_req_addr + 32'h3; // @[SimMem.scala 86:45]
  wire [31:0] _T_46 = _T_45 & 32'h3ffffff; // @[SimMem.scala 86:52]
  wire  _T_49 = 3'h3 == io_dcache_io_req_mtype; // @[Conditional.scala 37:30]
  wire [32:0] _T_50 = {{1'd0}, io_dcache_io_req_addr}; // @[SimMem.scala 91:47]
  wire [31:0] _T_52 = _T_50[31:0] & 32'h3ffffff; // @[SimMem.scala 91:54]
  wire [31:0] _T_71 = io_dcache_io_req_addr + 32'h4; // @[SimMem.scala 91:47]
  wire [31:0] _T_72 = _T_71 & 32'h3ffffff; // @[SimMem.scala 91:54]
  wire [31:0] _T_76 = io_dcache_io_req_addr + 32'h5; // @[SimMem.scala 91:47]
  wire [31:0] _T_77 = _T_76 & 32'h3ffffff; // @[SimMem.scala 91:54]
  wire [31:0] _T_81 = io_dcache_io_req_addr + 32'h6; // @[SimMem.scala 91:47]
  wire [31:0] _T_82 = _T_81 & 32'h3ffffff; // @[SimMem.scala 91:54]
  wire [31:0] _T_86 = io_dcache_io_req_addr + 32'h7; // @[SimMem.scala 91:47]
  wire [31:0] _T_87 = _T_86 & 32'h3ffffff; // @[SimMem.scala 91:54]
  wire  _T_90 = 3'h4 == io_dcache_io_req_mtype; // @[Conditional.scala 37:30]
  wire [31:0] _T_132 = io_dcache_io_req_addr + 32'h8; // @[SimMem.scala 97:47]
  wire [31:0] _T_133 = _T_132 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_137 = io_dcache_io_req_addr + 32'h9; // @[SimMem.scala 97:47]
  wire [31:0] _T_138 = _T_137 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_142 = io_dcache_io_req_addr + 32'ha; // @[SimMem.scala 97:47]
  wire [31:0] _T_143 = _T_142 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_147 = io_dcache_io_req_addr + 32'hb; // @[SimMem.scala 97:47]
  wire [31:0] _T_148 = _T_147 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_152 = io_dcache_io_req_addr + 32'hc; // @[SimMem.scala 97:47]
  wire [31:0] _T_153 = _T_152 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_157 = io_dcache_io_req_addr + 32'hd; // @[SimMem.scala 97:47]
  wire [31:0] _T_158 = _T_157 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_162 = io_dcache_io_req_addr + 32'he; // @[SimMem.scala 97:47]
  wire [31:0] _T_163 = _T_162 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_167 = io_dcache_io_req_addr + 32'hf; // @[SimMem.scala 97:47]
  wire [31:0] _T_168 = _T_167 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_172 = io_dcache_io_req_addr + 32'h10; // @[SimMem.scala 97:47]
  wire [31:0] _T_173 = _T_172 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_177 = io_dcache_io_req_addr + 32'h11; // @[SimMem.scala 97:47]
  wire [31:0] _T_178 = _T_177 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_182 = io_dcache_io_req_addr + 32'h12; // @[SimMem.scala 97:47]
  wire [31:0] _T_183 = _T_182 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_187 = io_dcache_io_req_addr + 32'h13; // @[SimMem.scala 97:47]
  wire [31:0] _T_188 = _T_187 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_192 = io_dcache_io_req_addr + 32'h14; // @[SimMem.scala 97:47]
  wire [31:0] _T_193 = _T_192 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_197 = io_dcache_io_req_addr + 32'h15; // @[SimMem.scala 97:47]
  wire [31:0] _T_198 = _T_197 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_202 = io_dcache_io_req_addr + 32'h16; // @[SimMem.scala 97:47]
  wire [31:0] _T_203 = _T_202 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_207 = io_dcache_io_req_addr + 32'h17; // @[SimMem.scala 97:47]
  wire [31:0] _T_208 = _T_207 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_212 = io_dcache_io_req_addr + 32'h18; // @[SimMem.scala 97:47]
  wire [31:0] _T_213 = _T_212 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_217 = io_dcache_io_req_addr + 32'h19; // @[SimMem.scala 97:47]
  wire [31:0] _T_218 = _T_217 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_222 = io_dcache_io_req_addr + 32'h1a; // @[SimMem.scala 97:47]
  wire [31:0] _T_223 = _T_222 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_227 = io_dcache_io_req_addr + 32'h1b; // @[SimMem.scala 97:47]
  wire [31:0] _T_228 = _T_227 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_232 = io_dcache_io_req_addr + 32'h1c; // @[SimMem.scala 97:47]
  wire [31:0] _T_233 = _T_232 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_237 = io_dcache_io_req_addr + 32'h1d; // @[SimMem.scala 97:47]
  wire [31:0] _T_238 = _T_237 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_242 = io_dcache_io_req_addr + 32'h1e; // @[SimMem.scala 97:47]
  wire [31:0] _T_243 = _T_242 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire [31:0] _T_247 = io_dcache_io_req_addr + 32'h1f; // @[SimMem.scala 97:47]
  wire [31:0] _T_248 = _T_247 & 32'h3ffffff; // @[SimMem.scala 97:54]
  wire  _GEN_122 = _T_49 ? 1'h0 : _T_90; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_200 = _T_30 ? 1'h0 : _T_49; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_219 = _T_30 ? 1'h0 : _GEN_122; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_293 = _T_21 ? 1'h0 : _T_30; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_304 = _T_21 ? 1'h0 : _GEN_200; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_323 = _T_21 ? 1'h0 : _GEN_219; // @[Conditional.scala 39:67 SimMem.scala 42:19]
  wire  _GEN_395 = _T_17 ? 1'h0 : _T_21; // @[Conditional.scala 40:58 SimMem.scala 42:19]
  wire  _GEN_402 = _T_17 ? 1'h0 : _GEN_293; // @[Conditional.scala 40:58 SimMem.scala 42:19]
  wire  _GEN_413 = _T_17 ? 1'h0 : _GEN_304; // @[Conditional.scala 40:58 SimMem.scala 42:19]
  wire  _GEN_432 = _T_17 ? 1'h0 : _GEN_323; // @[Conditional.scala 40:58 SimMem.scala 42:19]
  assign memory_icandidates_0_MPORT_addr = _icandidates_0_T_2[25:0];
  assign memory_icandidates_0_MPORT_data = memory[memory_icandidates_0_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_0_MPORT_addr = _dcandidates_0_T_3[25:0];
  assign memory_dcandidates_0_MPORT_data = memory[memory_dcandidates_0_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_1_MPORT_addr = _icandidates_1_T_2[25:0];
  assign memory_icandidates_1_MPORT_data = memory[memory_icandidates_1_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_1_MPORT_addr = _dcandidates_1_T_3[25:0];
  assign memory_dcandidates_1_MPORT_data = memory[memory_dcandidates_1_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_2_MPORT_addr = _icandidates_2_T_2[25:0];
  assign memory_icandidates_2_MPORT_data = memory[memory_icandidates_2_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_2_MPORT_addr = _dcandidates_2_T_3[25:0];
  assign memory_dcandidates_2_MPORT_data = memory[memory_dcandidates_2_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_3_MPORT_addr = _icandidates_3_T_2[25:0];
  assign memory_icandidates_3_MPORT_data = memory[memory_icandidates_3_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_3_MPORT_addr = _dcandidates_3_T_3[25:0];
  assign memory_dcandidates_3_MPORT_data = memory[memory_dcandidates_3_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_4_MPORT_addr = _icandidates_4_T_2[25:0];
  assign memory_icandidates_4_MPORT_data = memory[memory_icandidates_4_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_4_MPORT_addr = _dcandidates_4_T_3[25:0];
  assign memory_dcandidates_4_MPORT_data = memory[memory_dcandidates_4_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_5_MPORT_addr = _icandidates_5_T_2[25:0];
  assign memory_icandidates_5_MPORT_data = memory[memory_icandidates_5_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_5_MPORT_addr = _dcandidates_5_T_3[25:0];
  assign memory_dcandidates_5_MPORT_data = memory[memory_dcandidates_5_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_6_MPORT_addr = _icandidates_6_T_2[25:0];
  assign memory_icandidates_6_MPORT_data = memory[memory_icandidates_6_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_6_MPORT_addr = _dcandidates_6_T_3[25:0];
  assign memory_dcandidates_6_MPORT_data = memory[memory_dcandidates_6_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_7_MPORT_addr = _icandidates_7_T_2[25:0];
  assign memory_icandidates_7_MPORT_data = memory[memory_icandidates_7_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_7_MPORT_addr = _dcandidates_7_T_3[25:0];
  assign memory_dcandidates_7_MPORT_data = memory[memory_dcandidates_7_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_8_MPORT_addr = _icandidates_8_T_2[25:0];
  assign memory_icandidates_8_MPORT_data = memory[memory_icandidates_8_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_8_MPORT_addr = _dcandidates_8_T_3[25:0];
  assign memory_dcandidates_8_MPORT_data = memory[memory_dcandidates_8_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_9_MPORT_addr = _icandidates_9_T_2[25:0];
  assign memory_icandidates_9_MPORT_data = memory[memory_icandidates_9_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_9_MPORT_addr = _dcandidates_9_T_3[25:0];
  assign memory_dcandidates_9_MPORT_data = memory[memory_dcandidates_9_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_10_MPORT_addr = _icandidates_10_T_2[25:0];
  assign memory_icandidates_10_MPORT_data = memory[memory_icandidates_10_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_10_MPORT_addr = _dcandidates_10_T_3[25:0];
  assign memory_dcandidates_10_MPORT_data = memory[memory_dcandidates_10_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_11_MPORT_addr = _icandidates_11_T_2[25:0];
  assign memory_icandidates_11_MPORT_data = memory[memory_icandidates_11_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_11_MPORT_addr = _dcandidates_11_T_3[25:0];
  assign memory_dcandidates_11_MPORT_data = memory[memory_dcandidates_11_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_12_MPORT_addr = _icandidates_12_T_2[25:0];
  assign memory_icandidates_12_MPORT_data = memory[memory_icandidates_12_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_12_MPORT_addr = _dcandidates_12_T_3[25:0];
  assign memory_dcandidates_12_MPORT_data = memory[memory_dcandidates_12_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_13_MPORT_addr = _icandidates_13_T_2[25:0];
  assign memory_icandidates_13_MPORT_data = memory[memory_icandidates_13_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_13_MPORT_addr = _dcandidates_13_T_3[25:0];
  assign memory_dcandidates_13_MPORT_data = memory[memory_dcandidates_13_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_14_MPORT_addr = _icandidates_14_T_2[25:0];
  assign memory_icandidates_14_MPORT_data = memory[memory_icandidates_14_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_14_MPORT_addr = _dcandidates_14_T_3[25:0];
  assign memory_dcandidates_14_MPORT_data = memory[memory_dcandidates_14_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_15_MPORT_addr = _icandidates_15_T_2[25:0];
  assign memory_icandidates_15_MPORT_data = memory[memory_icandidates_15_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_15_MPORT_addr = _dcandidates_15_T_3[25:0];
  assign memory_dcandidates_15_MPORT_data = memory[memory_dcandidates_15_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_16_MPORT_addr = _icandidates_16_T_2[25:0];
  assign memory_icandidates_16_MPORT_data = memory[memory_icandidates_16_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_16_MPORT_addr = _dcandidates_16_T_3[25:0];
  assign memory_dcandidates_16_MPORT_data = memory[memory_dcandidates_16_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_17_MPORT_addr = _icandidates_17_T_2[25:0];
  assign memory_icandidates_17_MPORT_data = memory[memory_icandidates_17_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_17_MPORT_addr = _dcandidates_17_T_3[25:0];
  assign memory_dcandidates_17_MPORT_data = memory[memory_dcandidates_17_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_18_MPORT_addr = _icandidates_18_T_2[25:0];
  assign memory_icandidates_18_MPORT_data = memory[memory_icandidates_18_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_18_MPORT_addr = _dcandidates_18_T_3[25:0];
  assign memory_dcandidates_18_MPORT_data = memory[memory_dcandidates_18_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_19_MPORT_addr = _icandidates_19_T_2[25:0];
  assign memory_icandidates_19_MPORT_data = memory[memory_icandidates_19_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_19_MPORT_addr = _dcandidates_19_T_3[25:0];
  assign memory_dcandidates_19_MPORT_data = memory[memory_dcandidates_19_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_20_MPORT_addr = _icandidates_20_T_2[25:0];
  assign memory_icandidates_20_MPORT_data = memory[memory_icandidates_20_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_20_MPORT_addr = _dcandidates_20_T_3[25:0];
  assign memory_dcandidates_20_MPORT_data = memory[memory_dcandidates_20_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_21_MPORT_addr = _icandidates_21_T_2[25:0];
  assign memory_icandidates_21_MPORT_data = memory[memory_icandidates_21_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_21_MPORT_addr = _dcandidates_21_T_3[25:0];
  assign memory_dcandidates_21_MPORT_data = memory[memory_dcandidates_21_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_22_MPORT_addr = _icandidates_22_T_2[25:0];
  assign memory_icandidates_22_MPORT_data = memory[memory_icandidates_22_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_22_MPORT_addr = _dcandidates_22_T_3[25:0];
  assign memory_dcandidates_22_MPORT_data = memory[memory_dcandidates_22_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_23_MPORT_addr = _icandidates_23_T_2[25:0];
  assign memory_icandidates_23_MPORT_data = memory[memory_icandidates_23_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_23_MPORT_addr = _dcandidates_23_T_3[25:0];
  assign memory_dcandidates_23_MPORT_data = memory[memory_dcandidates_23_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_24_MPORT_addr = _icandidates_24_T_2[25:0];
  assign memory_icandidates_24_MPORT_data = memory[memory_icandidates_24_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_24_MPORT_addr = _dcandidates_24_T_3[25:0];
  assign memory_dcandidates_24_MPORT_data = memory[memory_dcandidates_24_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_25_MPORT_addr = _icandidates_25_T_2[25:0];
  assign memory_icandidates_25_MPORT_data = memory[memory_icandidates_25_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_25_MPORT_addr = _dcandidates_25_T_3[25:0];
  assign memory_dcandidates_25_MPORT_data = memory[memory_dcandidates_25_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_26_MPORT_addr = _icandidates_26_T_2[25:0];
  assign memory_icandidates_26_MPORT_data = memory[memory_icandidates_26_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_26_MPORT_addr = _dcandidates_26_T_3[25:0];
  assign memory_dcandidates_26_MPORT_data = memory[memory_dcandidates_26_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_27_MPORT_addr = _icandidates_27_T_2[25:0];
  assign memory_icandidates_27_MPORT_data = memory[memory_icandidates_27_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_27_MPORT_addr = _dcandidates_27_T_3[25:0];
  assign memory_dcandidates_27_MPORT_data = memory[memory_dcandidates_27_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_28_MPORT_addr = _icandidates_28_T_2[25:0];
  assign memory_icandidates_28_MPORT_data = memory[memory_icandidates_28_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_28_MPORT_addr = _dcandidates_28_T_3[25:0];
  assign memory_dcandidates_28_MPORT_data = memory[memory_dcandidates_28_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_29_MPORT_addr = _icandidates_29_T_2[25:0];
  assign memory_icandidates_29_MPORT_data = memory[memory_icandidates_29_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_29_MPORT_addr = _dcandidates_29_T_3[25:0];
  assign memory_dcandidates_29_MPORT_data = memory[memory_dcandidates_29_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_30_MPORT_addr = _icandidates_30_T_2[25:0];
  assign memory_icandidates_30_MPORT_data = memory[memory_icandidates_30_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_30_MPORT_addr = _dcandidates_30_T_3[25:0];
  assign memory_dcandidates_30_MPORT_data = memory[memory_dcandidates_30_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_icandidates_31_MPORT_addr = _icandidates_31_T_2[25:0];
  assign memory_icandidates_31_MPORT_data = memory[memory_icandidates_31_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_dcandidates_31_MPORT_addr = _dcandidates_31_T_3[25:0];
  assign memory_dcandidates_31_MPORT_data = memory[memory_dcandidates_31_MPORT_addr]; // @[SimMem.scala 42:19]
  assign memory_MPORT_data = io_dcache_io_req_data[7:0];
  assign memory_MPORT_addr = _T_18[25:0];
  assign memory_MPORT_mask = 1'h1;
  assign memory_MPORT_en = _T_16 & _T_17;
  assign memory_MPORT_1_data = io_dcache_io_req_data[7:0];
  assign memory_MPORT_1_addr = _T_18[25:0];
  assign memory_MPORT_1_mask = 1'h1;
  assign memory_MPORT_1_en = _T_16 & _GEN_395;
  assign memory_MPORT_2_data = io_dcache_io_req_data[15:8];
  assign memory_MPORT_2_addr = _T_27[25:0];
  assign memory_MPORT_2_mask = 1'h1;
  assign memory_MPORT_2_en = _T_16 & _GEN_395;
  assign memory_MPORT_3_data = io_dcache_io_req_data[7:0];
  assign memory_MPORT_3_addr = _T_18[25:0];
  assign memory_MPORT_3_mask = 1'h1;
  assign memory_MPORT_3_en = _T_16 & _GEN_402;
  assign memory_MPORT_4_data = io_dcache_io_req_data[15:8];
  assign memory_MPORT_4_addr = _T_27[25:0];
  assign memory_MPORT_4_mask = 1'h1;
  assign memory_MPORT_4_en = _T_16 & _GEN_402;
  assign memory_MPORT_5_data = io_dcache_io_req_data[23:16];
  assign memory_MPORT_5_addr = _T_41[25:0];
  assign memory_MPORT_5_mask = 1'h1;
  assign memory_MPORT_5_en = _T_16 & _GEN_402;
  assign memory_MPORT_6_data = io_dcache_io_req_data[31:24];
  assign memory_MPORT_6_addr = _T_46[25:0];
  assign memory_MPORT_6_mask = 1'h1;
  assign memory_MPORT_6_en = _T_16 & _GEN_402;
  assign memory_MPORT_7_data = io_dcache_io_req_data[7:0];
  assign memory_MPORT_7_addr = _T_52[25:0];
  assign memory_MPORT_7_mask = 1'h1;
  assign memory_MPORT_7_en = _T_16 & _GEN_413;
  assign memory_MPORT_8_data = io_dcache_io_req_data[15:8];
  assign memory_MPORT_8_addr = _T_27[25:0];
  assign memory_MPORT_8_mask = 1'h1;
  assign memory_MPORT_8_en = _T_16 & _GEN_413;
  assign memory_MPORT_9_data = io_dcache_io_req_data[23:16];
  assign memory_MPORT_9_addr = _T_41[25:0];
  assign memory_MPORT_9_mask = 1'h1;
  assign memory_MPORT_9_en = _T_16 & _GEN_413;
  assign memory_MPORT_10_data = io_dcache_io_req_data[31:24];
  assign memory_MPORT_10_addr = _T_46[25:0];
  assign memory_MPORT_10_mask = 1'h1;
  assign memory_MPORT_10_en = _T_16 & _GEN_413;
  assign memory_MPORT_11_data = io_dcache_io_req_data[39:32];
  assign memory_MPORT_11_addr = _T_72[25:0];
  assign memory_MPORT_11_mask = 1'h1;
  assign memory_MPORT_11_en = _T_16 & _GEN_413;
  assign memory_MPORT_12_data = io_dcache_io_req_data[47:40];
  assign memory_MPORT_12_addr = _T_77[25:0];
  assign memory_MPORT_12_mask = 1'h1;
  assign memory_MPORT_12_en = _T_16 & _GEN_413;
  assign memory_MPORT_13_data = io_dcache_io_req_data[55:48];
  assign memory_MPORT_13_addr = _T_82[25:0];
  assign memory_MPORT_13_mask = 1'h1;
  assign memory_MPORT_13_en = _T_16 & _GEN_413;
  assign memory_MPORT_14_data = io_dcache_io_req_data[63:56];
  assign memory_MPORT_14_addr = _T_87[25:0];
  assign memory_MPORT_14_mask = 1'h1;
  assign memory_MPORT_14_en = _T_16 & _GEN_413;
  assign memory_MPORT_15_data = io_dcache_io_req_data[7:0];
  assign memory_MPORT_15_addr = _T_52[25:0];
  assign memory_MPORT_15_mask = 1'h1;
  assign memory_MPORT_15_en = _T_16 & _GEN_432;
  assign memory_MPORT_16_data = io_dcache_io_req_data[15:8];
  assign memory_MPORT_16_addr = _T_27[25:0];
  assign memory_MPORT_16_mask = 1'h1;
  assign memory_MPORT_16_en = _T_16 & _GEN_432;
  assign memory_MPORT_17_data = io_dcache_io_req_data[23:16];
  assign memory_MPORT_17_addr = _T_41[25:0];
  assign memory_MPORT_17_mask = 1'h1;
  assign memory_MPORT_17_en = _T_16 & _GEN_432;
  assign memory_MPORT_18_data = io_dcache_io_req_data[31:24];
  assign memory_MPORT_18_addr = _T_46[25:0];
  assign memory_MPORT_18_mask = 1'h1;
  assign memory_MPORT_18_en = _T_16 & _GEN_432;
  assign memory_MPORT_19_data = io_dcache_io_req_data[39:32];
  assign memory_MPORT_19_addr = _T_72[25:0];
  assign memory_MPORT_19_mask = 1'h1;
  assign memory_MPORT_19_en = _T_16 & _GEN_432;
  assign memory_MPORT_20_data = io_dcache_io_req_data[47:40];
  assign memory_MPORT_20_addr = _T_77[25:0];
  assign memory_MPORT_20_mask = 1'h1;
  assign memory_MPORT_20_en = _T_16 & _GEN_432;
  assign memory_MPORT_21_data = io_dcache_io_req_data[55:48];
  assign memory_MPORT_21_addr = _T_82[25:0];
  assign memory_MPORT_21_mask = 1'h1;
  assign memory_MPORT_21_en = _T_16 & _GEN_432;
  assign memory_MPORT_22_data = io_dcache_io_req_data[63:56];
  assign memory_MPORT_22_addr = _T_87[25:0];
  assign memory_MPORT_22_mask = 1'h1;
  assign memory_MPORT_22_en = _T_16 & _GEN_432;
  assign memory_MPORT_23_data = io_dcache_io_req_data[71:64];
  assign memory_MPORT_23_addr = _T_133[25:0];
  assign memory_MPORT_23_mask = 1'h1;
  assign memory_MPORT_23_en = _T_16 & _GEN_432;
  assign memory_MPORT_24_data = io_dcache_io_req_data[79:72];
  assign memory_MPORT_24_addr = _T_138[25:0];
  assign memory_MPORT_24_mask = 1'h1;
  assign memory_MPORT_24_en = _T_16 & _GEN_432;
  assign memory_MPORT_25_data = io_dcache_io_req_data[87:80];
  assign memory_MPORT_25_addr = _T_143[25:0];
  assign memory_MPORT_25_mask = 1'h1;
  assign memory_MPORT_25_en = _T_16 & _GEN_432;
  assign memory_MPORT_26_data = io_dcache_io_req_data[95:88];
  assign memory_MPORT_26_addr = _T_148[25:0];
  assign memory_MPORT_26_mask = 1'h1;
  assign memory_MPORT_26_en = _T_16 & _GEN_432;
  assign memory_MPORT_27_data = io_dcache_io_req_data[103:96];
  assign memory_MPORT_27_addr = _T_153[25:0];
  assign memory_MPORT_27_mask = 1'h1;
  assign memory_MPORT_27_en = _T_16 & _GEN_432;
  assign memory_MPORT_28_data = io_dcache_io_req_data[111:104];
  assign memory_MPORT_28_addr = _T_158[25:0];
  assign memory_MPORT_28_mask = 1'h1;
  assign memory_MPORT_28_en = _T_16 & _GEN_432;
  assign memory_MPORT_29_data = io_dcache_io_req_data[119:112];
  assign memory_MPORT_29_addr = _T_163[25:0];
  assign memory_MPORT_29_mask = 1'h1;
  assign memory_MPORT_29_en = _T_16 & _GEN_432;
  assign memory_MPORT_30_data = io_dcache_io_req_data[127:120];
  assign memory_MPORT_30_addr = _T_168[25:0];
  assign memory_MPORT_30_mask = 1'h1;
  assign memory_MPORT_30_en = _T_16 & _GEN_432;
  assign memory_MPORT_31_data = io_dcache_io_req_data[135:128];
  assign memory_MPORT_31_addr = _T_173[25:0];
  assign memory_MPORT_31_mask = 1'h1;
  assign memory_MPORT_31_en = _T_16 & _GEN_432;
  assign memory_MPORT_32_data = io_dcache_io_req_data[143:136];
  assign memory_MPORT_32_addr = _T_178[25:0];
  assign memory_MPORT_32_mask = 1'h1;
  assign memory_MPORT_32_en = _T_16 & _GEN_432;
  assign memory_MPORT_33_data = io_dcache_io_req_data[151:144];
  assign memory_MPORT_33_addr = _T_183[25:0];
  assign memory_MPORT_33_mask = 1'h1;
  assign memory_MPORT_33_en = _T_16 & _GEN_432;
  assign memory_MPORT_34_data = io_dcache_io_req_data[159:152];
  assign memory_MPORT_34_addr = _T_188[25:0];
  assign memory_MPORT_34_mask = 1'h1;
  assign memory_MPORT_34_en = _T_16 & _GEN_432;
  assign memory_MPORT_35_data = io_dcache_io_req_data[167:160];
  assign memory_MPORT_35_addr = _T_193[25:0];
  assign memory_MPORT_35_mask = 1'h1;
  assign memory_MPORT_35_en = _T_16 & _GEN_432;
  assign memory_MPORT_36_data = io_dcache_io_req_data[175:168];
  assign memory_MPORT_36_addr = _T_198[25:0];
  assign memory_MPORT_36_mask = 1'h1;
  assign memory_MPORT_36_en = _T_16 & _GEN_432;
  assign memory_MPORT_37_data = io_dcache_io_req_data[183:176];
  assign memory_MPORT_37_addr = _T_203[25:0];
  assign memory_MPORT_37_mask = 1'h1;
  assign memory_MPORT_37_en = _T_16 & _GEN_432;
  assign memory_MPORT_38_data = io_dcache_io_req_data[191:184];
  assign memory_MPORT_38_addr = _T_208[25:0];
  assign memory_MPORT_38_mask = 1'h1;
  assign memory_MPORT_38_en = _T_16 & _GEN_432;
  assign memory_MPORT_39_data = io_dcache_io_req_data[199:192];
  assign memory_MPORT_39_addr = _T_213[25:0];
  assign memory_MPORT_39_mask = 1'h1;
  assign memory_MPORT_39_en = _T_16 & _GEN_432;
  assign memory_MPORT_40_data = io_dcache_io_req_data[207:200];
  assign memory_MPORT_40_addr = _T_218[25:0];
  assign memory_MPORT_40_mask = 1'h1;
  assign memory_MPORT_40_en = _T_16 & _GEN_432;
  assign memory_MPORT_41_data = io_dcache_io_req_data[215:208];
  assign memory_MPORT_41_addr = _T_223[25:0];
  assign memory_MPORT_41_mask = 1'h1;
  assign memory_MPORT_41_en = _T_16 & _GEN_432;
  assign memory_MPORT_42_data = io_dcache_io_req_data[223:216];
  assign memory_MPORT_42_addr = _T_228[25:0];
  assign memory_MPORT_42_mask = 1'h1;
  assign memory_MPORT_42_en = _T_16 & _GEN_432;
  assign memory_MPORT_43_data = io_dcache_io_req_data[231:224];
  assign memory_MPORT_43_addr = _T_233[25:0];
  assign memory_MPORT_43_mask = 1'h1;
  assign memory_MPORT_43_en = _T_16 & _GEN_432;
  assign memory_MPORT_44_data = io_dcache_io_req_data[239:232];
  assign memory_MPORT_44_addr = _T_238[25:0];
  assign memory_MPORT_44_mask = 1'h1;
  assign memory_MPORT_44_en = _T_16 & _GEN_432;
  assign memory_MPORT_45_data = io_dcache_io_req_data[247:240];
  assign memory_MPORT_45_addr = _T_243[25:0];
  assign memory_MPORT_45_mask = 1'h1;
  assign memory_MPORT_45_en = _T_16 & _GEN_432;
  assign memory_MPORT_46_data = io_dcache_io_req_data[255:248];
  assign memory_MPORT_46_addr = _T_248[25:0];
  assign memory_MPORT_46_mask = 1'h1;
  assign memory_MPORT_46_en = _T_16 & _GEN_432;
  assign io_icache_io_resp_valid = io_icache_io_resp_valid_REG; // @[SimMem.scala 63:27]
  assign io_icache_io_resp_data = io_icache_io_resp_data_REG; // @[SimMem.scala 64:27]
  assign io_dcache_io_resp_valid = io_dcache_io_resp_valid_REG; // @[SimMem.scala 65:27]
  assign io_dcache_io_resp_data = io_dcache_io_resp_data_REG; // @[SimMem.scala 66:27]
  always @(posedge clock) begin
    if(memory_MPORT_en & memory_MPORT_mask) begin
      memory[memory_MPORT_addr] <= memory_MPORT_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_1_en & memory_MPORT_1_mask) begin
      memory[memory_MPORT_1_addr] <= memory_MPORT_1_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_2_en & memory_MPORT_2_mask) begin
      memory[memory_MPORT_2_addr] <= memory_MPORT_2_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_3_en & memory_MPORT_3_mask) begin
      memory[memory_MPORT_3_addr] <= memory_MPORT_3_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_4_en & memory_MPORT_4_mask) begin
      memory[memory_MPORT_4_addr] <= memory_MPORT_4_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_5_en & memory_MPORT_5_mask) begin
      memory[memory_MPORT_5_addr] <= memory_MPORT_5_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_6_en & memory_MPORT_6_mask) begin
      memory[memory_MPORT_6_addr] <= memory_MPORT_6_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_7_en & memory_MPORT_7_mask) begin
      memory[memory_MPORT_7_addr] <= memory_MPORT_7_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_8_en & memory_MPORT_8_mask) begin
      memory[memory_MPORT_8_addr] <= memory_MPORT_8_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_9_en & memory_MPORT_9_mask) begin
      memory[memory_MPORT_9_addr] <= memory_MPORT_9_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_10_en & memory_MPORT_10_mask) begin
      memory[memory_MPORT_10_addr] <= memory_MPORT_10_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_11_en & memory_MPORT_11_mask) begin
      memory[memory_MPORT_11_addr] <= memory_MPORT_11_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_12_en & memory_MPORT_12_mask) begin
      memory[memory_MPORT_12_addr] <= memory_MPORT_12_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_13_en & memory_MPORT_13_mask) begin
      memory[memory_MPORT_13_addr] <= memory_MPORT_13_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_14_en & memory_MPORT_14_mask) begin
      memory[memory_MPORT_14_addr] <= memory_MPORT_14_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_15_en & memory_MPORT_15_mask) begin
      memory[memory_MPORT_15_addr] <= memory_MPORT_15_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_16_en & memory_MPORT_16_mask) begin
      memory[memory_MPORT_16_addr] <= memory_MPORT_16_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_17_en & memory_MPORT_17_mask) begin
      memory[memory_MPORT_17_addr] <= memory_MPORT_17_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_18_en & memory_MPORT_18_mask) begin
      memory[memory_MPORT_18_addr] <= memory_MPORT_18_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_19_en & memory_MPORT_19_mask) begin
      memory[memory_MPORT_19_addr] <= memory_MPORT_19_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_20_en & memory_MPORT_20_mask) begin
      memory[memory_MPORT_20_addr] <= memory_MPORT_20_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_21_en & memory_MPORT_21_mask) begin
      memory[memory_MPORT_21_addr] <= memory_MPORT_21_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_22_en & memory_MPORT_22_mask) begin
      memory[memory_MPORT_22_addr] <= memory_MPORT_22_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_23_en & memory_MPORT_23_mask) begin
      memory[memory_MPORT_23_addr] <= memory_MPORT_23_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_24_en & memory_MPORT_24_mask) begin
      memory[memory_MPORT_24_addr] <= memory_MPORT_24_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_25_en & memory_MPORT_25_mask) begin
      memory[memory_MPORT_25_addr] <= memory_MPORT_25_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_26_en & memory_MPORT_26_mask) begin
      memory[memory_MPORT_26_addr] <= memory_MPORT_26_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_27_en & memory_MPORT_27_mask) begin
      memory[memory_MPORT_27_addr] <= memory_MPORT_27_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_28_en & memory_MPORT_28_mask) begin
      memory[memory_MPORT_28_addr] <= memory_MPORT_28_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_29_en & memory_MPORT_29_mask) begin
      memory[memory_MPORT_29_addr] <= memory_MPORT_29_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_30_en & memory_MPORT_30_mask) begin
      memory[memory_MPORT_30_addr] <= memory_MPORT_30_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_31_en & memory_MPORT_31_mask) begin
      memory[memory_MPORT_31_addr] <= memory_MPORT_31_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_32_en & memory_MPORT_32_mask) begin
      memory[memory_MPORT_32_addr] <= memory_MPORT_32_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_33_en & memory_MPORT_33_mask) begin
      memory[memory_MPORT_33_addr] <= memory_MPORT_33_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_34_en & memory_MPORT_34_mask) begin
      memory[memory_MPORT_34_addr] <= memory_MPORT_34_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_35_en & memory_MPORT_35_mask) begin
      memory[memory_MPORT_35_addr] <= memory_MPORT_35_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_36_en & memory_MPORT_36_mask) begin
      memory[memory_MPORT_36_addr] <= memory_MPORT_36_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_37_en & memory_MPORT_37_mask) begin
      memory[memory_MPORT_37_addr] <= memory_MPORT_37_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_38_en & memory_MPORT_38_mask) begin
      memory[memory_MPORT_38_addr] <= memory_MPORT_38_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_39_en & memory_MPORT_39_mask) begin
      memory[memory_MPORT_39_addr] <= memory_MPORT_39_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_40_en & memory_MPORT_40_mask) begin
      memory[memory_MPORT_40_addr] <= memory_MPORT_40_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_41_en & memory_MPORT_41_mask) begin
      memory[memory_MPORT_41_addr] <= memory_MPORT_41_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_42_en & memory_MPORT_42_mask) begin
      memory[memory_MPORT_42_addr] <= memory_MPORT_42_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_43_en & memory_MPORT_43_mask) begin
      memory[memory_MPORT_43_addr] <= memory_MPORT_43_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_44_en & memory_MPORT_44_mask) begin
      memory[memory_MPORT_44_addr] <= memory_MPORT_44_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_45_en & memory_MPORT_45_mask) begin
      memory[memory_MPORT_45_addr] <= memory_MPORT_45_data; // @[SimMem.scala 42:19]
    end
    if(memory_MPORT_46_en & memory_MPORT_46_mask) begin
      memory[memory_MPORT_46_addr] <= memory_MPORT_46_data; // @[SimMem.scala 42:19]
    end
    io_icache_io_resp_valid_REG <= io_icache_io_req_valid; // @[SimMem.scala 63:37]
    io_icache_io_resp_data_REG <= {io_icache_io_resp_data_hi,io_icache_io_resp_data_lo}; // @[SimMem.scala 64:50]
    io_dcache_io_resp_valid_REG <= io_dcache_io_req_valid; // @[SimMem.scala 65:37]
    io_dcache_io_resp_data_REG <= {io_dcache_io_resp_data_hi,io_dcache_io_resp_data_lo}; // @[SimMem.scala 66:50]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_dcache_io_req_valid & _T_6 & ~reset) begin
          $fwrite(32'h80000002,"%c",io_dcache_io_req_data[7:0]); // @[SimMem.scala 30:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_icache_io_req_valid & _T_10 & _T_9) begin
          $fwrite(32'h80000002,"icache is accessing %x, ram overflow\n",io_icache_io_req_addr); // @[SimMem.scala 36:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
  integer initvar;
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_icache_io_resp_valid_REG = _RAND_0[0:0];
  _RAND_1 = {8{`RANDOM}};
  io_icache_io_resp_data_REG = _RAND_1[255:0];
  _RAND_2 = {1{`RANDOM}};
  io_dcache_io_resp_valid_REG = _RAND_2[0:0];
  _RAND_3 = {8{`RANDOM}};
  io_dcache_io_resp_data_REG = _RAND_3[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
  $readmemh("testfile.hex", memory);
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TileForVerilator(
  input         clock,
  input         reset,
  output [63:0] io_difftest_gprs_0,
  output [63:0] io_difftest_gprs_1,
  output [63:0] io_difftest_gprs_2,
  output [63:0] io_difftest_gprs_3,
  output [63:0] io_difftest_gprs_4,
  output [63:0] io_difftest_gprs_5,
  output [63:0] io_difftest_gprs_6,
  output [63:0] io_difftest_gprs_7,
  output [63:0] io_difftest_gprs_8,
  output [63:0] io_difftest_gprs_9,
  output [63:0] io_difftest_gprs_10,
  output [63:0] io_difftest_gprs_11,
  output [63:0] io_difftest_gprs_12,
  output [63:0] io_difftest_gprs_13,
  output [63:0] io_difftest_gprs_14,
  output [63:0] io_difftest_gprs_15,
  output [63:0] io_difftest_gprs_16,
  output [63:0] io_difftest_gprs_17,
  output [63:0] io_difftest_gprs_18,
  output [63:0] io_difftest_gprs_19,
  output [63:0] io_difftest_gprs_20,
  output [63:0] io_difftest_gprs_21,
  output [63:0] io_difftest_gprs_22,
  output [63:0] io_difftest_gprs_23,
  output [63:0] io_difftest_gprs_24,
  output [63:0] io_difftest_gprs_25,
  output [63:0] io_difftest_gprs_26,
  output [63:0] io_difftest_gprs_27,
  output [63:0] io_difftest_gprs_28,
  output [63:0] io_difftest_gprs_29,
  output [63:0] io_difftest_gprs_30,
  output [63:0] io_difftest_gprs_31,
  output        io_difftest_valids_0,
  output        io_difftest_valids_1,
  output        io_difftest_valids_2,
  output [63:0] io_difftest_pcs_0,
  output [63:0] io_difftest_pcs_1,
  output [63:0] io_difftest_pcs_2,
  output [1:0]  io_difftest_orders_0,
  output [1:0]  io_difftest_orders_1,
  output [1:0]  io_difftest_orders_2,
  output [31:0] io_difftest_insts_0,
  output [31:0] io_difftest_insts_1,
  output [31:0] io_difftest_insts_2,
  output [63:0] io_difftest_csrs_mstatus,
  output [63:0] io_difftest_csrs_sstatus,
  output [63:0] io_difftest_csrs_mepc,
  output [63:0] io_difftest_csrs_sepc,
  output [63:0] io_difftest_csrs_mtval,
  output [63:0] io_difftest_csrs_stval,
  output [63:0] io_difftest_csrs_mtvec,
  output [63:0] io_difftest_csrs_stvec,
  output [63:0] io_difftest_csrs_mcause,
  output [63:0] io_difftest_csrs_scause,
  output [63:0] io_difftest_csrs_satp,
  output [63:0] io_difftest_csrs_mip,
  output [63:0] io_difftest_csrs_mie,
  output [63:0] io_difftest_csrs_mscratch,
  output [63:0] io_difftest_csrs_sscratch,
  output [63:0] io_difftest_csrs_mideleg,
  output [63:0] io_difftest_csrs_medeleg,
  output        io_difftest_int,
  input         io_difftest_sync,
  input  [4:0]  io_difftest_saddr,
  input  [31:0] io_difftest_sval,
  output        io_difftest_finish,
  output        io_difftest_mmio_0,
  output        io_difftest_mmio_1,
  output        io_difftest_mmio_2,
  output        io_difftest_print_0,
  output        io_difftest_print_1,
  output        io_difftest_print_2,
  output [1:0]  io_difftest_mode,
  output [63:0] io_difftest_counter,
  output [63:0] io_difftest_common,
  output [63:0] io_difftest_dstall,
  output [63:0] io_difftest_istall,
  output [63:0] io_difftest_mduStall,
  output [63:0] io_difftest_instret
);
  wire  core_clock; // @[Tile.scala 103:20]
  wire  core_reset; // @[Tile.scala 103:20]
  wire [31:0] core_io_icache_req_bits_addr; // @[Tile.scala 103:20]
  wire [2:0] core_io_icache_req_bits_mtype; // @[Tile.scala 103:20]
  wire  core_io_icache_resp_valid; // @[Tile.scala 103:20]
  wire [31:0] core_io_icache_resp_bits_rdata_0; // @[Tile.scala 103:20]
  wire [31:0] core_io_icache_resp_bits_rdata_1; // @[Tile.scala 103:20]
  wire  core_io_icache_resp_bits_respn; // @[Tile.scala 103:20]
  wire  core_io_dcache_req_valid; // @[Tile.scala 103:20]
  wire [31:0] core_io_dcache_req_bits_addr; // @[Tile.scala 103:20]
  wire [63:0] core_io_dcache_req_bits_wdata; // @[Tile.scala 103:20]
  wire  core_io_dcache_req_bits_wen; // @[Tile.scala 103:20]
  wire [2:0] core_io_dcache_req_bits_mtype; // @[Tile.scala 103:20]
  wire  core_io_dcache_resp_valid; // @[Tile.scala 103:20]
  wire [31:0] core_io_dcache_resp_bits_rdata_0; // @[Tile.scala 103:20]
  wire [31:0] core_io_dcache_resp_bits_rdata_1; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mstatus; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_sstatus; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mepc; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_sepc; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mtval; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_stval; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mtvec; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_stvec; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mcause; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_scause; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_satp; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mip; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mie; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mscratch; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_sscratch; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_mideleg; // @[Tile.scala 103:20]
  wire [63:0] core_csrs_medeleg; // @[Tile.scala 103:20]
  wire [63:0] core_istall; // @[Tile.scala 103:20]
  wire  core__WIRE_4_0; // @[Tile.scala 103:20]
  wire  core__WIRE_4_1; // @[Tile.scala 103:20]
  wire  core__WIRE_4_2; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_1_0; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_1_1; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_1_2; // @[Tile.scala 103:20]
  wire [4:0] core_difftest_saddr; // @[Tile.scala 103:20]
  wire [1:0] core_current_mode; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__0; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__1; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__2; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__3; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__4; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__5; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__6; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__7; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__8; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__9; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__10; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__11; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__12; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__13; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__14; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__15; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__16; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__17; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__18; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__19; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__20; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__21; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__22; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__23; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__24; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__25; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__26; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__27; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__28; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__29; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__30; // @[Tile.scala 103:20]
  wire [63:0] core__WIRE__31; // @[Tile.scala 103:20]
  wire [63:0] core_dstall; // @[Tile.scala 103:20]
  wire  core__WIRE_0_0; // @[Tile.scala 103:20]
  wire  core__WIRE_0_1; // @[Tile.scala 103:20]
  wire  core__WIRE_0_2; // @[Tile.scala 103:20]
  wire [63:0] core_counter; // @[Tile.scala 103:20]
  wire [31:0] core_difftest_sval; // @[Tile.scala 103:20]
  wire [63:0] core_mduStall; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_3_0; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_3_1; // @[Tile.scala 103:20]
  wire [31:0] core__WIRE_3_2; // @[Tile.scala 103:20]
  wire [63:0] core_common; // @[Tile.scala 103:20]
  wire  core__WIRE_5_0; // @[Tile.scala 103:20]
  wire  core__WIRE_5_1; // @[Tile.scala 103:20]
  wire  core__WIRE_5_2; // @[Tile.scala 103:20]
  wire [63:0] core_instret; // @[Tile.scala 103:20]
  wire [1:0] core__WIRE_2_0; // @[Tile.scala 103:20]
  wire [1:0] core__WIRE_2_1; // @[Tile.scala 103:20]
  wire [1:0] core__WIRE_2_2; // @[Tile.scala 103:20]
  wire  core_REG_0; // @[Tile.scala 103:20]
  wire  core_difftest_sync; // @[Tile.scala 103:20]
  wire  core_wbInsts_0_ysyx_debug; // @[Tile.scala 103:20]
  wire  icache_clock; // @[Tile.scala 104:22]
  wire  icache_reset; // @[Tile.scala 104:22]
  wire [31:0] icache_io_cpu_req_bits_addr; // @[Tile.scala 104:22]
  wire [2:0] icache_io_cpu_req_bits_mtype; // @[Tile.scala 104:22]
  wire  icache_io_cpu_resp_valid; // @[Tile.scala 104:22]
  wire [31:0] icache_io_cpu_resp_bits_rdata_0; // @[Tile.scala 104:22]
  wire [31:0] icache_io_cpu_resp_bits_rdata_1; // @[Tile.scala 104:22]
  wire  icache_io_cpu_resp_bits_respn; // @[Tile.scala 104:22]
  wire  icache_io_bar_req_valid; // @[Tile.scala 104:22]
  wire [31:0] icache_io_bar_req_addr; // @[Tile.scala 104:22]
  wire  icache_io_bar_resp_valid; // @[Tile.scala 104:22]
  wire [255:0] icache_io_bar_resp_data; // @[Tile.scala 104:22]
  wire  dcache_clock; // @[Tile.scala 105:22]
  wire  dcache_reset; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_cpu_req_valid; // @[Tile.scala 105:22]
  wire [31:0] dcache_io_dcache_cpu_req_bits_addr; // @[Tile.scala 105:22]
  wire [63:0] dcache_io_dcache_cpu_req_bits_wdata; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_cpu_req_bits_wen; // @[Tile.scala 105:22]
  wire [2:0] dcache_io_dcache_cpu_req_bits_mtype; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_cpu_resp_valid; // @[Tile.scala 105:22]
  wire [31:0] dcache_io_dcache_cpu_resp_bits_rdata_0; // @[Tile.scala 105:22]
  wire [31:0] dcache_io_dcache_cpu_resp_bits_rdata_1; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_bar_req_valid; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_bar_req_wen; // @[Tile.scala 105:22]
  wire [31:0] dcache_io_dcache_bar_req_addr; // @[Tile.scala 105:22]
  wire [255:0] dcache_io_dcache_bar_req_data; // @[Tile.scala 105:22]
  wire [2:0] dcache_io_dcache_bar_req_mtype; // @[Tile.scala 105:22]
  wire  dcache_io_dcache_bar_resp_valid; // @[Tile.scala 105:22]
  wire [255:0] dcache_io_dcache_bar_resp_data; // @[Tile.scala 105:22]
  wire  mem_clock; // @[Tile.scala 106:19]
  wire  mem_reset; // @[Tile.scala 106:19]
  wire  mem_io_icache_io_req_valid; // @[Tile.scala 106:19]
  wire [31:0] mem_io_icache_io_req_addr; // @[Tile.scala 106:19]
  wire  mem_io_icache_io_resp_valid; // @[Tile.scala 106:19]
  wire [255:0] mem_io_icache_io_resp_data; // @[Tile.scala 106:19]
  wire  mem_io_dcache_io_req_valid; // @[Tile.scala 106:19]
  wire  mem_io_dcache_io_req_wen; // @[Tile.scala 106:19]
  wire [31:0] mem_io_dcache_io_req_addr; // @[Tile.scala 106:19]
  wire [255:0] mem_io_dcache_io_req_data; // @[Tile.scala 106:19]
  wire [2:0] mem_io_dcache_io_req_mtype; // @[Tile.scala 106:19]
  wire  mem_io_dcache_io_resp_valid; // @[Tile.scala 106:19]
  wire [255:0] mem_io_dcache_io_resp_data; // @[Tile.scala 106:19]
  wire  difftest__sync = io_difftest_sync;
  wire [31:0] difftest__sval = io_difftest_sval;
  wire [4:0] difftest__saddr = io_difftest_saddr;
  wire [31:0] difftestPCs_0 = core__WIRE_1_0;
  wire [31:0] difftestPCs_1 = core__WIRE_1_1;
  wire [31:0] difftestPCs_2 = core__WIRE_1_2;
  Core core ( // @[Tile.scala 103:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_icache_req_bits_addr(core_io_icache_req_bits_addr),
    .io_icache_req_bits_mtype(core_io_icache_req_bits_mtype),
    .io_icache_resp_valid(core_io_icache_resp_valid),
    .io_icache_resp_bits_rdata_0(core_io_icache_resp_bits_rdata_0),
    .io_icache_resp_bits_rdata_1(core_io_icache_resp_bits_rdata_1),
    .io_icache_resp_bits_respn(core_io_icache_resp_bits_respn),
    .io_dcache_req_valid(core_io_dcache_req_valid),
    .io_dcache_req_bits_addr(core_io_dcache_req_bits_addr),
    .io_dcache_req_bits_wdata(core_io_dcache_req_bits_wdata),
    .io_dcache_req_bits_wen(core_io_dcache_req_bits_wen),
    .io_dcache_req_bits_mtype(core_io_dcache_req_bits_mtype),
    .io_dcache_resp_valid(core_io_dcache_resp_valid),
    .io_dcache_resp_bits_rdata_0(core_io_dcache_resp_bits_rdata_0),
    .io_dcache_resp_bits_rdata_1(core_io_dcache_resp_bits_rdata_1),
    .csrs_mstatus(core_csrs_mstatus),
    .csrs_sstatus(core_csrs_sstatus),
    .csrs_mepc(core_csrs_mepc),
    .csrs_sepc(core_csrs_sepc),
    .csrs_mtval(core_csrs_mtval),
    .csrs_stval(core_csrs_stval),
    .csrs_mtvec(core_csrs_mtvec),
    .csrs_stvec(core_csrs_stvec),
    .csrs_mcause(core_csrs_mcause),
    .csrs_scause(core_csrs_scause),
    .csrs_satp(core_csrs_satp),
    .csrs_mip(core_csrs_mip),
    .csrs_mie(core_csrs_mie),
    .csrs_mscratch(core_csrs_mscratch),
    .csrs_sscratch(core_csrs_sscratch),
    .csrs_mideleg(core_csrs_mideleg),
    .csrs_medeleg(core_csrs_medeleg),
    .istall(core_istall),
    ._WIRE_4_0(core__WIRE_4_0),
    ._WIRE_4_1(core__WIRE_4_1),
    ._WIRE_4_2(core__WIRE_4_2),
    ._WIRE_1_0(core__WIRE_1_0),
    ._WIRE_1_1(core__WIRE_1_1),
    ._WIRE_1_2(core__WIRE_1_2),
    .difftest_saddr(core_difftest_saddr),
    .current_mode(core_current_mode),
    ._WIRE__0(core__WIRE__0),
    ._WIRE__1(core__WIRE__1),
    ._WIRE__2(core__WIRE__2),
    ._WIRE__3(core__WIRE__3),
    ._WIRE__4(core__WIRE__4),
    ._WIRE__5(core__WIRE__5),
    ._WIRE__6(core__WIRE__6),
    ._WIRE__7(core__WIRE__7),
    ._WIRE__8(core__WIRE__8),
    ._WIRE__9(core__WIRE__9),
    ._WIRE__10(core__WIRE__10),
    ._WIRE__11(core__WIRE__11),
    ._WIRE__12(core__WIRE__12),
    ._WIRE__13(core__WIRE__13),
    ._WIRE__14(core__WIRE__14),
    ._WIRE__15(core__WIRE__15),
    ._WIRE__16(core__WIRE__16),
    ._WIRE__17(core__WIRE__17),
    ._WIRE__18(core__WIRE__18),
    ._WIRE__19(core__WIRE__19),
    ._WIRE__20(core__WIRE__20),
    ._WIRE__21(core__WIRE__21),
    ._WIRE__22(core__WIRE__22),
    ._WIRE__23(core__WIRE__23),
    ._WIRE__24(core__WIRE__24),
    ._WIRE__25(core__WIRE__25),
    ._WIRE__26(core__WIRE__26),
    ._WIRE__27(core__WIRE__27),
    ._WIRE__28(core__WIRE__28),
    ._WIRE__29(core__WIRE__29),
    ._WIRE__30(core__WIRE__30),
    ._WIRE__31(core__WIRE__31),
    .dstall(core_dstall),
    ._WIRE_0_0(core__WIRE_0_0),
    ._WIRE_0_1(core__WIRE_0_1),
    ._WIRE_0_2(core__WIRE_0_2),
    .counter(core_counter),
    .difftest_sval(core_difftest_sval),
    .mduStall(core_mduStall),
    ._WIRE_3_0(core__WIRE_3_0),
    ._WIRE_3_1(core__WIRE_3_1),
    ._WIRE_3_2(core__WIRE_3_2),
    .common(core_common),
    ._WIRE_5_0(core__WIRE_5_0),
    ._WIRE_5_1(core__WIRE_5_1),
    ._WIRE_5_2(core__WIRE_5_2),
    .instret(core_instret),
    ._WIRE_2_0(core__WIRE_2_0),
    ._WIRE_2_1(core__WIRE_2_1),
    ._WIRE_2_2(core__WIRE_2_2),
    .REG_0(core_REG_0),
    .difftest_sync(core_difftest_sync),
    .wbInsts_0_ysyx_debug(core_wbInsts_0_ysyx_debug)
  );
  ICache icache ( // @[Tile.scala 104:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_cpu_req_bits_addr(icache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_mtype(icache_io_cpu_req_bits_mtype),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_rdata_0(icache_io_cpu_resp_bits_rdata_0),
    .io_cpu_resp_bits_rdata_1(icache_io_cpu_resp_bits_rdata_1),
    .io_cpu_resp_bits_respn(icache_io_cpu_resp_bits_respn),
    .io_bar_req_valid(icache_io_bar_req_valid),
    .io_bar_req_addr(icache_io_bar_req_addr),
    .io_bar_resp_valid(icache_io_bar_resp_valid),
    .io_bar_resp_data(icache_io_bar_resp_data)
  );
  DcacheDPFilter dcache ( // @[Tile.scala 105:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dcache_cpu_req_valid(dcache_io_dcache_cpu_req_valid),
    .io_dcache_cpu_req_bits_addr(dcache_io_dcache_cpu_req_bits_addr),
    .io_dcache_cpu_req_bits_wdata(dcache_io_dcache_cpu_req_bits_wdata),
    .io_dcache_cpu_req_bits_wen(dcache_io_dcache_cpu_req_bits_wen),
    .io_dcache_cpu_req_bits_mtype(dcache_io_dcache_cpu_req_bits_mtype),
    .io_dcache_cpu_resp_valid(dcache_io_dcache_cpu_resp_valid),
    .io_dcache_cpu_resp_bits_rdata_0(dcache_io_dcache_cpu_resp_bits_rdata_0),
    .io_dcache_cpu_resp_bits_rdata_1(dcache_io_dcache_cpu_resp_bits_rdata_1),
    .io_dcache_bar_req_valid(dcache_io_dcache_bar_req_valid),
    .io_dcache_bar_req_wen(dcache_io_dcache_bar_req_wen),
    .io_dcache_bar_req_addr(dcache_io_dcache_bar_req_addr),
    .io_dcache_bar_req_data(dcache_io_dcache_bar_req_data),
    .io_dcache_bar_req_mtype(dcache_io_dcache_bar_req_mtype),
    .io_dcache_bar_resp_valid(dcache_io_dcache_bar_resp_valid),
    .io_dcache_bar_resp_data(dcache_io_dcache_bar_resp_data)
  );
  SimMem mem ( // @[Tile.scala 106:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_icache_io_req_valid(mem_io_icache_io_req_valid),
    .io_icache_io_req_addr(mem_io_icache_io_req_addr),
    .io_icache_io_resp_valid(mem_io_icache_io_resp_valid),
    .io_icache_io_resp_data(mem_io_icache_io_resp_data),
    .io_dcache_io_req_valid(mem_io_dcache_io_req_valid),
    .io_dcache_io_req_wen(mem_io_dcache_io_req_wen),
    .io_dcache_io_req_addr(mem_io_dcache_io_req_addr),
    .io_dcache_io_req_data(mem_io_dcache_io_req_data),
    .io_dcache_io_req_mtype(mem_io_dcache_io_req_mtype),
    .io_dcache_io_resp_valid(mem_io_dcache_io_resp_valid),
    .io_dcache_io_resp_data(mem_io_dcache_io_resp_data)
  );
  assign io_difftest_gprs_0 = core__WIRE__0; // @[Tile.scala 141:15]
  assign io_difftest_gprs_1 = core__WIRE__1; // @[Tile.scala 141:15]
  assign io_difftest_gprs_2 = core__WIRE__2; // @[Tile.scala 141:15]
  assign io_difftest_gprs_3 = core__WIRE__3; // @[Tile.scala 141:15]
  assign io_difftest_gprs_4 = core__WIRE__4; // @[Tile.scala 141:15]
  assign io_difftest_gprs_5 = core__WIRE__5; // @[Tile.scala 141:15]
  assign io_difftest_gprs_6 = core__WIRE__6; // @[Tile.scala 141:15]
  assign io_difftest_gprs_7 = core__WIRE__7; // @[Tile.scala 141:15]
  assign io_difftest_gprs_8 = core__WIRE__8; // @[Tile.scala 141:15]
  assign io_difftest_gprs_9 = core__WIRE__9; // @[Tile.scala 141:15]
  assign io_difftest_gprs_10 = core__WIRE__10; // @[Tile.scala 141:15]
  assign io_difftest_gprs_11 = core__WIRE__11; // @[Tile.scala 141:15]
  assign io_difftest_gprs_12 = core__WIRE__12; // @[Tile.scala 141:15]
  assign io_difftest_gprs_13 = core__WIRE__13; // @[Tile.scala 141:15]
  assign io_difftest_gprs_14 = core__WIRE__14; // @[Tile.scala 141:15]
  assign io_difftest_gprs_15 = core__WIRE__15; // @[Tile.scala 141:15]
  assign io_difftest_gprs_16 = core__WIRE__16; // @[Tile.scala 141:15]
  assign io_difftest_gprs_17 = core__WIRE__17; // @[Tile.scala 141:15]
  assign io_difftest_gprs_18 = core__WIRE__18; // @[Tile.scala 141:15]
  assign io_difftest_gprs_19 = core__WIRE__19; // @[Tile.scala 141:15]
  assign io_difftest_gprs_20 = core__WIRE__20; // @[Tile.scala 141:15]
  assign io_difftest_gprs_21 = core__WIRE__21; // @[Tile.scala 141:15]
  assign io_difftest_gprs_22 = core__WIRE__22; // @[Tile.scala 141:15]
  assign io_difftest_gprs_23 = core__WIRE__23; // @[Tile.scala 141:15]
  assign io_difftest_gprs_24 = core__WIRE__24; // @[Tile.scala 141:15]
  assign io_difftest_gprs_25 = core__WIRE__25; // @[Tile.scala 141:15]
  assign io_difftest_gprs_26 = core__WIRE__26; // @[Tile.scala 141:15]
  assign io_difftest_gprs_27 = core__WIRE__27; // @[Tile.scala 141:15]
  assign io_difftest_gprs_28 = core__WIRE__28; // @[Tile.scala 141:15]
  assign io_difftest_gprs_29 = core__WIRE__29; // @[Tile.scala 141:15]
  assign io_difftest_gprs_30 = core__WIRE__30; // @[Tile.scala 141:15]
  assign io_difftest_gprs_31 = core__WIRE__31; // @[Tile.scala 141:15]
  assign io_difftest_valids_0 = core__WIRE_0_0; // @[Tile.scala 141:15]
  assign io_difftest_valids_1 = core__WIRE_0_1; // @[Tile.scala 141:15]
  assign io_difftest_valids_2 = core__WIRE_0_2; // @[Tile.scala 141:15]
  assign io_difftest_pcs_0 = {{32'd0}, difftestPCs_0}; // @[Tile.scala 141:15]
  assign io_difftest_pcs_1 = {{32'd0}, difftestPCs_1}; // @[Tile.scala 141:15]
  assign io_difftest_pcs_2 = {{32'd0}, difftestPCs_2}; // @[Tile.scala 141:15]
  assign io_difftest_orders_0 = core__WIRE_2_0; // @[Tile.scala 141:15]
  assign io_difftest_orders_1 = core__WIRE_2_1; // @[Tile.scala 141:15]
  assign io_difftest_orders_2 = core__WIRE_2_2; // @[Tile.scala 141:15]
  assign io_difftest_insts_0 = core__WIRE_3_0; // @[Tile.scala 141:15]
  assign io_difftest_insts_1 = core__WIRE_3_1; // @[Tile.scala 141:15]
  assign io_difftest_insts_2 = core__WIRE_3_2; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mstatus = core_csrs_mstatus; // @[Tile.scala 141:15]
  assign io_difftest_csrs_sstatus = core_csrs_sstatus; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mepc = core_csrs_mepc; // @[Tile.scala 141:15]
  assign io_difftest_csrs_sepc = core_csrs_sepc; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mtval = core_csrs_mtval; // @[Tile.scala 141:15]
  assign io_difftest_csrs_stval = core_csrs_stval; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mtvec = core_csrs_mtvec; // @[Tile.scala 141:15]
  assign io_difftest_csrs_stvec = core_csrs_stvec; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mcause = core_csrs_mcause; // @[Tile.scala 141:15]
  assign io_difftest_csrs_scause = core_csrs_scause; // @[Tile.scala 141:15]
  assign io_difftest_csrs_satp = core_csrs_satp; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mip = core_csrs_mip; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mie = core_csrs_mie; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mscratch = core_csrs_mscratch; // @[Tile.scala 141:15]
  assign io_difftest_csrs_sscratch = core_csrs_sscratch; // @[Tile.scala 141:15]
  assign io_difftest_csrs_mideleg = core_csrs_mideleg; // @[Tile.scala 141:15]
  assign io_difftest_csrs_medeleg = core_csrs_medeleg; // @[Tile.scala 141:15]
  assign io_difftest_int = core_REG_0; // @[Tile.scala 141:15]
  assign io_difftest_finish = core_wbInsts_0_ysyx_debug; // @[Tile.scala 141:15]
  assign io_difftest_mmio_0 = core__WIRE_4_0; // @[Tile.scala 141:15]
  assign io_difftest_mmio_1 = core__WIRE_4_1; // @[Tile.scala 141:15]
  assign io_difftest_mmio_2 = core__WIRE_4_2; // @[Tile.scala 141:15]
  assign io_difftest_print_0 = core__WIRE_5_0; // @[Tile.scala 141:15]
  assign io_difftest_print_1 = core__WIRE_5_1; // @[Tile.scala 141:15]
  assign io_difftest_print_2 = core__WIRE_5_2; // @[Tile.scala 141:15]
  assign io_difftest_mode = core_current_mode; // @[Tile.scala 141:15]
  assign io_difftest_counter = core_counter; // @[Tile.scala 141:15]
  assign io_difftest_common = core_common; // @[Tile.scala 141:15]
  assign io_difftest_dstall = core_dstall; // @[Tile.scala 141:15]
  assign io_difftest_istall = core_istall; // @[Tile.scala 141:15]
  assign io_difftest_mduStall = core_mduStall; // @[Tile.scala 141:15]
  assign io_difftest_instret = core_instret; // @[Tile.scala 141:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_icache_resp_valid = icache_io_cpu_resp_valid; // @[Tile.scala 111:18]
  assign core_io_icache_resp_bits_rdata_0 = icache_io_cpu_resp_bits_rdata_0; // @[Tile.scala 111:18]
  assign core_io_icache_resp_bits_rdata_1 = icache_io_cpu_resp_bits_rdata_1; // @[Tile.scala 111:18]
  assign core_io_icache_resp_bits_respn = icache_io_cpu_resp_bits_respn; // @[Tile.scala 111:18]
  assign core_io_dcache_resp_valid = dcache_io_dcache_cpu_resp_valid; // @[Tile.scala 112:18]
  assign core_io_dcache_resp_bits_rdata_0 = dcache_io_dcache_cpu_resp_bits_rdata_0; // @[Tile.scala 112:18]
  assign core_io_dcache_resp_bits_rdata_1 = dcache_io_dcache_cpu_resp_bits_rdata_1; // @[Tile.scala 112:18]
  assign core_difftest_saddr = difftest__saddr;
  assign core_difftest_sval = difftest__sval;
  assign core_difftest_sync = difftest__sync;
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_cpu_req_bits_addr = core_io_icache_req_bits_addr; // @[Tile.scala 111:18]
  assign icache_io_cpu_req_bits_mtype = core_io_icache_req_bits_mtype; // @[Tile.scala 111:18]
  assign icache_io_bar_resp_valid = mem_io_icache_io_resp_valid; // @[Tile.scala 113:20]
  assign icache_io_bar_resp_data = mem_io_icache_io_resp_data; // @[Tile.scala 113:20]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dcache_cpu_req_valid = core_io_dcache_req_valid; // @[Tile.scala 112:18]
  assign dcache_io_dcache_cpu_req_bits_addr = core_io_dcache_req_bits_addr; // @[Tile.scala 112:18]
  assign dcache_io_dcache_cpu_req_bits_wdata = core_io_dcache_req_bits_wdata; // @[Tile.scala 112:18]
  assign dcache_io_dcache_cpu_req_bits_wen = core_io_dcache_req_bits_wen; // @[Tile.scala 112:18]
  assign dcache_io_dcache_cpu_req_bits_mtype = core_io_dcache_req_bits_mtype; // @[Tile.scala 112:18]
  assign dcache_io_dcache_bar_resp_valid = mem_io_dcache_io_resp_valid; // @[Tile.scala 114:20]
  assign dcache_io_dcache_bar_resp_data = mem_io_dcache_io_resp_data; // @[Tile.scala 114:20]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_icache_io_req_valid = icache_io_bar_req_valid; // @[Tile.scala 113:20]
  assign mem_io_icache_io_req_addr = icache_io_bar_req_addr; // @[Tile.scala 113:20]
  assign mem_io_dcache_io_req_valid = dcache_io_dcache_bar_req_valid; // @[Tile.scala 114:20]
  assign mem_io_dcache_io_req_wen = dcache_io_dcache_bar_req_wen; // @[Tile.scala 114:20]
  assign mem_io_dcache_io_req_addr = dcache_io_dcache_bar_req_addr; // @[Tile.scala 114:20]
  assign mem_io_dcache_io_req_data = dcache_io_dcache_bar_req_data; // @[Tile.scala 114:20]
  assign mem_io_dcache_io_req_mtype = dcache_io_dcache_bar_req_mtype; // @[Tile.scala 114:20]
endmodule
